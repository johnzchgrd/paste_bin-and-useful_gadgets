
//////////////////////////////////////////////////////////////////////////////////
// Company       : 
// Engineer      : Johnzchgrd
// 
// Create Date   : 2020-08-07 18:21:52
// Design Name   : 
// File Name     : lcd_ctrl.v
// Project Name  : 
// Target Devices: Tang Nano(GW1N-LV1QN48C5/I4)
// Tool Versions : 
// Description   : a generic LCD display controller.
// 
// Dependencies  : -
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module lcd_ctrl (
  input        clk  , // <=25.2MHz, tested 10.2MHz~24MHz, recommended <20MHz for more stable display
  input        rst  ,
  output       DE   , // data enable
  output       hsync,
  output       vsync,
  output [9:0] h_cnt,
  output [9:0] v_cnt
);

/* timing parameters */
parameter pixel_height = 'd272;
parameter pixel_width  = 'd480;
/* copied from szg's lecture */
// see note in the bottom of this file.
localparam v_p = 'd2         ;
localparam v_q = 'd33        ;
localparam v_r = pixel_height;
localparam v_s = 'd10        ;

localparam h_b = 'd77       ;
localparam h_c = 'd53       ;
localparam h_d = pixel_width;
localparam h_e = 'd24       ;

/* extreme situation also works... no idea why...
localparam v_p = 'd1         ;
localparam v_q = 'd0         ;
localparam v_r = pixel_height;
localparam v_s = 'd1         ;

localparam h_b = 'd1        ;
localparam h_c = 'd0        ;
localparam h_d = pixel_width;
localparam h_e = 'd1        ;
*/

localparam v_p_q     = v_p     + v_q;
localparam v_p_q_r   = v_p_q   + v_r;
localparam v_p_q_r_s = v_p_q_r + v_s;
localparam h_b_c     = h_b     + h_c;
localparam h_b_c_d   = h_b_c   + h_d;
localparam h_b_c_d_e = h_b_c_d + h_e;

/* nets definitions */
reg  [9:0] pcnt_h ; // pixel counts
reg  [9:0] pcnt_v ;
wire       h_valid;
wire       v_valid;


always@(posedge clk or posedge rst) begin
  if(rst) begin
    pcnt_v <= 'd1;
    pcnt_h <= 'd1;
  end else begin
    pcnt_h <= pcnt_h == h_b_c_d_e ? 'd1 : pcnt_h + 'd1;
    pcnt_v <= pcnt_h == h_b_c_d_e ?
      (pcnt_v == v_p_q_r_s ? 'd1 : pcnt_v + 'd1) :
      pcnt_v;
  end
end

assign h_valid = (pcnt_h > h_b_c && pcnt_h <= h_b_c_d) ? 1'b1 :
                 1'b0;
assign v_valid = (pcnt_v > v_p_q && pcnt_v <= v_p_q_r) ? 1'b1 : 
                 1'b0; 
assign DE = h_valid & v_valid;

/* generate VSYNC & HSYNC */

assign hsync = (pcnt_h <= h_b ? 1'b1 : 1'b0);
assign vsync = (pcnt_v <= v_p ? 1'b1 : 1'b0);

assign h_cnt = h_valid ? pcnt_h - h_b_c : 'd0;
assign v_cnt = v_valid ? pcnt_v - v_p_q : 'd0;
 
endmodule


// note for meaning of those "strange" identifiers:
/* use "http://tool.chinaz.com/tools/imgtobase/" to decode
data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAAtIAAAFqCAYAAAA3G70vAAAAAXNSR0IArs4c6QAAAARnQU1BAACxjwv8YQUAAAAJcEhZcwAADsMAAA7DAcdvqGQAAOYiSURBVHhe7N0HmGRVtf/949V7r1lREAVRAck5KjnnIEjOknPOWXIOA0OQKIOkIeecc85JgglFVEC9il7/17fe+uw6e7qm6Zmuqq7urula3+epp7tOnbjPDr+99tprf6JSpQiCIAiCIAiCoCn+o/wbBEEQBEEQBEEThJAOgiAIgiAIghYIIR0EQRAEQRAELRBCOgiCIAiCIAhaIIR0EARBEARBELRACOkgCIIgCIIgaIEQ0kEQBEEQBEHQAiGkgyAIgiAIgqAFYkGWIAiCNvH//X//X/HnP/+5+OUvf1luCYKgk/j85z9fTDvttMV//ud/lluCYGCEkA6CBvl//+//FS+++GLxX//1X8Xss89ebu1eiMY//elPxZNPPlmsssoq5dbu5o9//GNx0kknFe+//37x2c9+ttw6cVTB//rXv4q//vWvxRRTTFFu7R/p/9FHHxX//ve/iy996Uvl1v75v//7v+Ivf/lL8YUvfCHl5UaR/z/44INiyimnLLf0z1Dfo3T88MMPW7pHf7/4xS+WW/tHevzP//xPEmbN3qPO1te+9rVyS/8M5B7lq8997nPFpz/96XJr//zv//5vSv9m7tE7do/yc7P3+Pe//z3dX7P32GyZcS0stdRSxTrrrJP+73Z+85vfFK+99lqx3HLLlVuCZgkhHQQNouK+7777iv/+7/8ullxyyXJr96JR//Wvf13cdNNNxU477VRu7W7eeOONYuWVVy7WXHPNYo455ii3Thyi8c033yxuvvnmYs899yy39g/R8thjjyXB43qN8oc//KG45pprihVWWCFZ5hrFuz7//POLww47rNzSP3/729+Kxx9/PAnONdZYo9zaP7///e+L66+/Pt3jd77znXJr/xgJGDNmTHHIIYeUW/rHvblH6bn66quXW/vnd7/7XXpnyy+/fPHtb3+73No/b731VnH55ZcXBx54YLmlfwjGJ554ovjnP/9ZrLrqquXW/nnnnXeKG2+8sVhkkUWKOeecs9zaPz//+c9THtlvv/3KLf0jH7pHYlUZaJR333031auME42WGbz66qup7tl7773LLf2jo3vPPfcUU001VXHOOeeUW7ubV155pXjkkUeKrbbaqtwSNA0hHQRB//zrX/+qPPvss5WXXnqp3NLd/Pvf/6689957lVtuuaXcElQFSGWuueaq3HHHHeWW/pGv7r333spyyy1XbmmMDz74oDJ69OjKQQcdVG5pjKqQq6y33nqVqugptzSGvD/33HOX3xrj/fffr5x++umVqrAttzTG66+/Xtlggw0qTz31VLmlMZ588snK/PPPX35rjKq4qpx22mmVww8/vNzSGFUBUtl4440rTz/9dLmlMaqipbLQQguV3xpDORs1alTlqKOOKrc0xgsvvFBZd911K1XBX25pjPvvv7+y+OKLl98aoyqIK6ecckrlmGOOKbc0RlUQV3bbbbfKrbfeWm5pjLvvvruy9NJLl98ao9rRquyxxx6V7bbbrtwSVDvIlTvvvLP8FrRCTDYMggZhgWU9YdELahiSZYUNalTr1GSRYzkMgqCz4H6izuJeE9Qw2vH222+X34JWCCEdBA1CJHHv8Alq6ZH9IoMedLh8giDoLHKdFeWzB65lUYcPjBDSQdAgn/zkJ5O/5jTTTFNu6W4+8YlPpAlkc889d7klkCZ86BudaBgEwdDxqU99Kk1gbWZS40jnq1/9alO+6cHHCSEdBA3CiiEigEk1QQ0uDCZdBTVYvFh4cnSAIAg6B9ZoI4rKaFCDNdrk3qB1Qkh3GMTas88+W5x55pnllu5FAR89enSaUd8JeDfvvfdemvkd1ESjdxT+deNDRIf7TxB0HupwdVZ0dHvgIx1x7wdGCOkWISKIKmGWen9+/OMfF7feemu5Z+Mo5M8880wKL9VsaB6Wwfp7OProo1Ov+9FHHy33GH5UXkIP1d9n/hx++OHFHXfcUe5Ze54LL7ywOPbYY1Oc4k6Aa4dwYd/61rfKLd0NNwbxYuedd95ySxCuHUHQuXDt4I6mjAY1Jp988mKuueYqvwWtEEJ6AGg0fW677bbirrvuSoX0P/7jP4qXXnqpOPLII1sS044n2BqF+BaDlhC9++670z34ENEEfafFyvRsZkyfcMIJqSOS04xVU5qNHTs27Sdd/eZvJ6ED5RP0IA8G4xN5JAg6kyib4yM9og4fGCGkW4TAs+rTAQccUMw///zF9773vXHWVUHshQTLorBRCEpO/80sCmAImYh+6KGHknDO97DPPvuk81lEoVOwJOsSSyxR7LXXXskisMUWW4y7X9v+8Y9/FCeeeGLa1+9rr7128eUvfzl97wRUNnzJIvxdDRVwhL8bH2kSrh1B0JnkKEMR/q6HCH83cEJItxkNqeVfCe16F4BsOT700EPT56ijjip/qf3GLzpvb3Qym0rhueeeK66++upi5513Hm+JT7OSDzrooGK77bZL392XGMhE93XXXZfcR6644opx2/N9cQlx/2DVvvfee9P2vD9UQlbLuuyyy9IKWPk4q2i1AsE/9dRTp/8nm2yy9Lce9/jb3/42XeeYY45J1yHg6r8ju4PYLh3b7VvtPr/+9a83tWzuSEYet/TwDDPMUG4JpIkOY0QFCILOw4got6tmlnQf6XDPm2666cpvQSuEkG4DhDBf5Cw4+QHvuuuuxfrrrz/u91/84hdJiCrIhOGll16ahGgW0WefffY4l477778//e0PQpdfMReIvtbJV1mss8466X/WXhZrgje7oWj0WVh/8pOfpGu7F0ve+u7crNyWfPUbK5tjbSOunYsrxpVXXpmOu+WWW5qywBO93E6kmQ9L9CyzzDLB5V6lGVcQLiFENZzDcb7737K7nsdz6bQcf/zxLYv7vnBeAin863qQN4jpoAcdLp8gCDoPdVaUzx5ogZjTMTAiN7UJBZOFmIWUhZfLB2EI21lwf/azn6X/iVRDvybSEagENoGW3UIadWcgYH/zm98kgVd/jHOyOmeRyjpLUKpAfOabb77iwAMPLNZcc83igQceSMI53xfB7TtBesYZZxT33Xdf+o0V+vXXX0/COQsFBXCmmWYq9t9//2KRRRYpHnvssfIO+sc9Oz5Xan/729/SNd56661yjx7s+41vfKPYcsstyy1FEm977rln+j9brI877rh0fH4OPuPtnKgoHcxuluZBLd0NCxoVCWpIE2Xb8HEQBJ2FOlydxfAS1Hj//ffTvK6gdUJItwFCkI80Vwr+zcTbyy+/XP5aK7yvvvpqclsgHInmTTfdtNhwww2T6GXNXWWVVdK+fl988cXT//1BYJqBnAV1Pe5JmDbi8n/+53/SNbfeeut0/nqBzzXjK1/5Str+mc98plhjjTWSO4jfXnzxxSTQ/fb5z3++OPjgg4vFFlusWHjhhVOkBiKaH7P7MDzUDL19pFmiDYm7X2nVDJ5fZcAfXHqwxM8666xJ4H/zm98s9xo40lR6uEbQY6HXyQl60EGUl4Mg6CzU4eosZTSowRo95ZRTlt+CVggh3UYIOJZoopMVOPsaQwEmPLNwtJ+QM0Qgt49WUBkQ8Cy5rMgZjfiqq65abLPNNkmwEsYTEpTEEL/f+vsillnWnH+FFVYY95sJjFaFajfuQUFeb731kvjnTtIKOgJZnOvU+F/6tgvvUFpNMcUU5ZbuxntTCU8//fTllkCahI90EHQmjELhIz0+jGDCugatE0K6jRBalkved999k1sBH2JiOluBWapzXGfuB9lnWqSOMWPGpH0Jv+effz75A/e3KItjF1100WLllVcuLrjgguKss84qf2kMx88444zJKn377benbUQ59w1igFX32muvTW4hWfAPVkxnQ22XXHJJuqepppqq3NpDtgYT+CzsLPkmE3LhcJy/JgHmcH9+l9btXHUvXDvGJ1w7Pk527TAZNgiCzkK7G64d42M01+hz0DohpFtEg0nsioKRBTLhTOQRthtssEFx2mmnJR9l7gorrbRSEtMm6dnGP9o2FmOW3qeffjptP+KII8b5PROVruGYvkRytuSywPIfPv3008f5RfsQlfyhuSLweTahUSNPtBPHLM6E+LLLLpsmSTrGBD0C2nlZtIV6s93v/K6XWmqpNCHxqaeeSi4YRKwJiDoO+bvJiNKid9QM4tZv0kNFVj/Z0Pmvv/76YqeddioWXHDBJIzdr+vfeeedyUrNEswCf+6556bzZ1HvOVjcd9lllxTBxPn4qhO9ztVupHvQQ6THx4k0CYJgUkBdFfXVwAghPQBkPkJ4tdVWS+I5+10ZNiLquBd89atfTdZdw9++m5RHIHNDWHfdddMxjjf5z762b7bZZkk8E7IZQrLeVSTjXKzgzr399tun7z6uSVzyE2bJZdEVYs51vv3tb6dj3T9XBdtWXHHFdJxhL37P7kvMZ64e9vdMQuQQpoatf/CDH6SoJI7x25JLLjnuu2uxYBPAvfEb95B83ny/hpeIab7S2QfZfjvuuGOx0EILpeNMMDQZc7bZZkvptPTSS6djdESkL79z/zuf3x2Xw+q1A/cQrh3jE64d46NMKXsR2SUIOg9tg3YkXDt60M5+5zvfKb8FLVEJOpp//vOflUMPPbRyyimnVD788MNya+fyf//3f5WnnnqqUhW4lSuvvLLcOjLwLm699dbKPffcU27pbv79739XfvGLX1ROO+20ckvw+uuvV2adddbKjTfeWG7pn3/961+Ve++9t7LccsuVWxrjgw8+qIwePbpS7USXWxrjrbfeqqy33nqVaue83NIYzz77bKXaaS+/Ncb7779fOf300yuHHHJIuaUxpOMGG2yQ6pJmePLJJyvzzz9/+a0x/vjHP6Y8fPjhh5dbGuOVV16pbLzxxpWnn3663NIYjzzySKXayS+/NcZ7771XGTVqVOWoo44qtzTGCy+8UFl33XUrN998c7mlMe6///7K4osvXn5rjHfffTe1U8ccc0y5pTFeffXVym677Zbq1ma4++67K0svvXT5rTHk/W233bayxRZblFuCl156qXLOOeeU34JWCIv0JAALF+tqfYi7ToZVjtWay8hIolpekktKrFpXQ3rwORS6MOjBaAx/+iAIOgt1lrLZzknokzrq8JjTMTBCSHc4hoi5XvANnhQwdCY0HheLSUX4N4pnMwQ2zTTTlFu6Gx0mLjlci4Ia2d2Ly0sQBJ0Fl0WuDBFVpwcupQIeBK0TQjoIGoQVg596o0u4dwOs8yayBjWyld7E2iAIOgvWaHWWMhrUsHiUoAZB64SQDoIGIaSJRrGug5poVAlbjj3ogYgO958g6DzU4eqs6Oj2IBxgq2tZBDVCSAdBg3DtELg+XDtqZNcOrjxBjXDtCILOhWuHOiui6vQw+eSTF3POOWf5LWiFENJB0ASssMH4RJoEQRBMmkT9PXBCSAddicrDTGU+z41+Pvjgg+Ktt95Kw2B9/d5tnw8//DC5ulgVq6/fu/HDf97qoLFyWhB0Hnyk1fvN1v0j+fPb3/62eOmll/r8rRs/6nALwjXDJ6qCIrojQddB6Fii/dlnny239I9K2GqJhgfzojbdjKqDf90bb7xRzD///OXW7kZ6WKV09OjRxWKLLVZunTgmPmnIrAp6wgknlFv7R9jBu+66K3Xwtthii3Jr/1g2/7zzzivWW2+9YqaZZiq39g9feCuyOrZRpMfDDz+cFkiyaFOjWLb4vvvuS2E/p5pqqnJr/3i2m266abzFrPqDz6zOoDrBIlSNYq7Egw8+mO7xG9/4Rrm1f6wqe/vtt6fVaBuF8JNHdNIazVewMqw8YtGkZiI/vfDCC8X5559fjBo1qtzSP/LhPffck+5xww03LLf2z69//evixhtvLBZYYIGmVqJVd1988cXFySefXG7pH2lvxWGLhTXzrkcyf/rTn1K6RPSlGhbrkQ8tTNcoIaSDrsRkMJX3yy+/XG7pH4LH8u2EdPhJ1ybuWBL/7bffLuaZZ55ya3dDRBBmlrpvdMVHVTAryK9+9atirrnmKrf2j/xotr1r8t1vFNYWoyrysFBgjUK4v/baa011mkzqIqaF2MoQXNdee20636qrrjounTwHsa6zaqVY5H2lzzLLLDPB9CEYf/azn6X8+LWvfS2dl0CzkmxfsDzdcccd6fwbbbRRU+nQCsTKddddl6x/GSu4Wp2VfypR/uijjyaxO+WUU5Z79M+7775bXHnllUnIr7POOuXW8ZGu0vorX/lKuaV/pI880ky5dh3vQb3wrW99q9zaP8qLDpD7a+YejYgpM80IQM912223Fffff39apTao5U3pH37SNazboZ5ZZZVVyi39E0I6CBqExUolLAapJdW7HRZ6ja2G3FL0Qc2SevnllxcrrbRSWlI/GB/Cj0WQSxABVC+kbfMbMXz66acn8Xfvvfcm66EJYhq4bbfd9mMCiAhwnHPnNHes8uo8fUFQsWaOHTs2va+pp566/GVwIFYuvPDC4vrrr0/3+M1vfjMJfZZ6ZYeQb0VI69gfd9xxSYgbYQsmjvf++OOPJ7GvjAZF8fzzz6dytttuu5VbgmYJH+kgaBARGSwyo1EPeiJUhGWnB6MVLKIRFeDjsP7qdBGQ3Bp23XXXcSKalfzVV18dL54t6+att96aLK0s/DqwDz30UPlrDYKZOwF3mj322KM49NBDi+23375fC7NybGh/qMqyyAiGihdddNFi0003Tfe58cYbF6+88krxyCOPFFNMMUWx+uqrNyWi4bgVVlih/Bb0h8hL3nnU4T3ozKmzgtb55I+rlP8HQTARDN6wlgltFhVPLT0M50qTGWaYodza3XC34IbArzeHwJNOLGD/8R/da7cwekEo87nlhsLdQ7pkFwAim+WZZZhVnzj8+c9/nvydd9xxx5SWXADsk90+wLfznHPOKb7//e+P82n83Oc+l4ZmiVLnJ7bvvvvu4tJLL02+v0QtFwKi3faFF144XeeJJ55I741YJ+AJ92eeeSb97/51AriC2cc1n3zyySRk+S+ziHNx8lyXXXZZuuZ3v/vddD8Z1lCCn0XahwXe9e3HnSULaqNeV1999Ti/bZZm17CqKteaM888s3juuefSc3KZcV3Pteaaa6Y0Zmnn9iAdu90FLQ+46/TDe5SmOrpRh9dQrqRJjKC1Tlikg6BB8mRDw6lBrZEiHDTqQQ2+98RWFooEjWHTBx54oNyjO2Fx5v9sIg+Byw2D2wUxqePx1FNPFbPMMsu40Q0dEmmY4/7qhLAmEs71EJj8ZGecccZySw0WZ/7Rrku8EsfOSYieccYZ6br18F0+++yzU6eQG8Y111yTIvQQoybd+U255wryk5/8JIlwIttESp1J1zjxxBPTd/fomL5wvjFjxhSHHXZYcdFFFyWhT8hLDwLc9eUZLiA33HBDmmBIWCP7Q8O9EPP2z0gv6cjdyn3kfbsZ74mPPcu/+tu7knZRh/egEyufBa0TQjoIGoRVg5Uqhu1rSA9C5/Of/3y5JSD4WE9ZJFkyjznmmOKkk05K4ppFshs/xB6LF/FK3HLrEFWDCCZAuXDw8eX20AoE9oTyoOs/9thjKToJd4rNNtssRZnhF5ph1c1zHpzHjH0+zNxDRJLwP4G/9dZbJ7FPnHEf4c/sXKzIfL2998UXXzy5bOhw14vc3ig3zrXzzjsX8803XzrO9SabbLIUTWWHHXZI36XNfvvtlyZastBncey5TJhjjc4QidJR/eTcBDp0IOrfRzd9pI8OyxFHHJGizehI8bWPOrwHedHoRtA6MdkwCBpEBAKCSEU822yzlVu7F+4KrHfEUEzcqUFAcz9gAWNRJNg02mussUbXDp0SoWuttVayuOp88Xc2QZBFlUWWEBaizf+EKYsudw7pddRRRyWXDB2UW265JVn2hRbMEJf77rtvEprOmyGipD0XDtE8/L788sunc7Moc0Uy2dFEP/fBIk3c33zzzekdEl5EN9cI98CvefbZZ09uEyJkcC9xX6zW9mXBFgXoqquuSsKd0OYuUj+JkaXYtZdddtn0qYd1m5clyzfXEa4aP/rRj9L/3Eb8ZZk+6KCDxkXn0AEQ9cM9eEaTGbmnSCN+r1xouLvwSfdbN6JjId10bLw3IRjlA9FIvM+gNrrx+uuvfyxPBo0TFukgaBDCUQNtKDqowZWh9zB5N8P6p3PByiPWOH9csFcId9aNH5ZVll4TC/kBc0GQb6QTQcvVo7c/MXGdfZwJYmXO8HPvWNT24U/NFSJbmblz+D93YnxMSIThfe+od6fG+8oTFN1bbxeSoYT4I4h/8IMfpA77WWedlVxCWKuJ40022SRZqXuH5/JcBLTt0lungFXcs/X1XrrhIx10wowk6hTxizYSEnV4D8qLkY+gdcIiHQQNooHl76phXmqppcqt3YuORV5MwRB1UIttS9RZNEN+sagIQcddoJkFOEYi8grrLZ9nwoa/9O677z4uggJLMOshl4Uc/o51X/xlImhi4e9OOeWU5IPNyszqzVrLVYTvNGs3q67v8iwrtQgZLMqG/bfbbrskPlm2iX0uEqy69nc+FnCuF97pueeem67Pws1f2vncE79nVm3nyP7JLMz5ndeHv5t33nmLrbbaalzcXsKZJdqCPNw6uIqwZhPLJjTyvXaPrOAszzoiOmlEIrcQ/tgs89xBdGqlm7xHWB955JHjOgjdCFcOE1z5zOuEcfFhnfbeWPODIo2y6uByXQpaI6J2BEGD6HPqvWv4Y8Z3LT24u2i0I2pHDRZPs+BZUokdQmzWWWdNDbnh+W6GtVTkCS4OhC63g94rArJEE5LyE6FtP9Yywpv7UG/LNQhFw/R5sRPXyavkEd+s1qyTBCsRzZ/Zd0PaedTAvo4jUll+dZR95x/tO/Hs/bk/ot4xOtQsxuoC7927ti+RRiR7tuw+wApKwHk252IRd1+QX1jAszh2HJcQos9zu659iWbP7zk8l/9dRwfFX+fN5VBngviX97oZ1mjvUMdpjjnmSHlKnRWRl3pQf8u/EbWjdcIiHQQNwlKl564BtSxwt0MwEC9CePHnDIo0ZGzFPBO9BnuRjyAImoOrCwss4TihVS+7DaMZ5rlssMEG5ZagWcJHOggahHAMH+ke9MFZM4TlCmoYTmdBlS5BEHQWBLT6O+rwHoyy1i+EFDRPCOkgaBDDuoamu32Rg4zhY0PkZsAHNQzFG+6PldOCoPMwmqj+5kYT1OA+lf31g9YIIR0EDZItsGFt7IEFlv9nUMOoBZ9Xlq8gCDoL5TPq8PGJOnzghJAOggZRCXNjiFBBNXQsVMB87IIa/OhNpouGKQg6DxMN1d/hytADNxexyIPWCSEdBA1iBrhZ+dwZgpprB1eGmFTXg5i9IiwYQg6CoLPgnqf+jjq8BxFMekfPCZojhHQQNAHh6BPU0DAJ2RXU0Nmy3C5BHQRBZ6F86uRGHd6DUIqxRPjACCEdBA2SXTtiWLBGdu2wvGxQg2vH22+/Ha4dQdCBhGvHx+HaYTGjoHVCSAdBg+QoFRGRoYb0YN3pvdJcN8MSbdGNcO0Igs7DCJr6O+rwHiw8FIvTDIwQ0kHQICphvmRR6dQgpA0J9rXaXLdimHTaaadNfodBEHQWyqf6O+rwHnQqYlXDgRFCOggaREgzy/xazjeouXZYUvn5558vtwTCalk5zQpqQRB0Flyv1N+Whw9qfPDBB8VLL71UfgtaIYR0EDQJARn0EOkxPpEeQdC5RPkcH+kRaTIwQkgHQYOY8c0fOIYFe+DCEK4dPYRrRxB0LuYwhGvH+HDtUGcFrRNCOggaRK/9z3/+c3JnCGpwZYgZ8D1w//njH/8YK6cFQQeifKq/RaoIavzjH/9IdVbQOiGkg6BBCOl//vOf6RPU0DCFP3APQiT+7W9/iyXCg6ADyXV4dHR7EBJQnRW0ziQjpP/0pz8VRx11VMdMElAgxYs99thjk5WyUzCZ4tJLLy3uvPPOcsvgYp3+Bx54oDjvvPPKLe1BRXfZZZcVd999d7ll+AnXjo8Trh3jw7XjO9/5Trh2BEEHksNTRh3eQ7h2DJxPVAXhgL3Mf/WrXxUXXXRR+a0WJuzAAw9M1pkjjzyy3FrbvuOOOxZf/vKXyy2NQ0ifccYZxeabb15861vfKrcOD5JMUPd99tmnuOqqq9IsfY1nb4jMyy+/PAluDexqq62Wen4zzzxzS2nQH3qWN9xwQ3HQQQcVK6+8cnHSSSeVvwwenvGhhx5Ki3Jsu+225daBw2ogbVV4yy+/fLm1fehw3HPPPcXPf/7zckv/yM+GBBdbbLFi6aWXLrd2L9LjF7/4RepExRKzNZTB3//+98Xkk0+e4rMGQdA5aK/U4dpwZTQoio8++qiYbLLJiq222ipptJGCUUHa9P77729q1JRWm2WWWYoll1yy3NI/bRHSQoJpTIlGPZtFFlmk+PGPf5we5NBDDy1uu+22lHk32mijYtddd00vrVNR0K655ppi3XXXLbd8HEnGL3SvvfYqrr322j6FtGd/8MEHixNOOKGYb7750jbLkj7++OPFqFGj+hTeA0Uj7n4OOeSQYpVVVhkSId0uWKBvvvnm4oc//GG5ZXDhF3bFFVcUzz77bLmlf9yj97fGGmukfN3tyG86USrgVVddtdza3chXOpXqQYv3BEHQOajDrU6rDQ8rbA2j/NKDMXQkLVRDPN90001pZLuZd/1f//VfxYILLliss8465Zb+aYuQBgHK4rrMMsskgZkhKHfaaaf0sjxUJ8PCJiYusc9dYWJ4LhZNoqovIa3A7r777umlnHrqqSl9WIsvuOCCYvTo0YMipMHirROgRzWpCGnpLg0JMkJ1KHBNoxzNLOWsYHLlmWqqqYoTTzyx3Nq9sOrfd999xd57711cd9115dbuRn565plnillnnbX46le/Wm4NgqAT0NFlpVT/K6NBkXQMd1CfKaecstw66WMC5dixY4s33ngjabpG4cL5+c9/vqn6e1iEtEs+8sgj6QXCcMIBBxyQ/pfBWQr1jDRIftt+++2TRduL3mGHHdJvt956a/q9Hv5P+++/f7pmdqmQKHw411tvvbSP+zz++OOL1VdfPRUoFkk+U1tvvXWyrp122mnJkrzbbrsVP/jBD9JvZ599djrWvcw///zJ1aA/Ic014Uc/+lEaNjnuuOOSsHUMoTjTTDOloPCEtfubccYZi7XWWisNk+s9cWfYbLPNilNOOSVZlt3nc889lzK5+4TnYOl3/+7LOdZee+1xQtp31l3DGpYr3mabbVK6SZMrr7yymH322VMQ9gUWWCC5Kdju2rC/0YOpp546XefRRx8tXnvttfR+zz333PS79OOiwirJH1sF5XqGtXv7S+tMuMYcc8yRjudTnv2NPadnY6VnTT/44IPTvu5vzJgxxbzzzpvuUZ5hSTj//PPTOd2D9yMt3eMLL7yQntVznnzyyema8qL31S7cN9HILcdIQ7dDSEtzZe6pp54qt3Y3OlvqEfl2JDVKQTAS0NElrOgMZTQoki6jNUaikOYeSjccfvjh5dbBoa2TDYmdu+66qzjiiCPGfUwQrBe89nnxxReTVZYIIzh/+tOfFkcffXTK3Ib3DZvzrfa7xprlUEIcdthhxYcffpj2e/jhh9PvLL9PP/10+o0Y9Nstt9ySzuN3BcdvxDnBdfrppyfXB+d3H/n3V155JQldq/y4R9d1vHMR1q7z5JNPpudpZHIhUU/YPvbYY+neWTK90IUXXji5trgX4tT5/A/Xc9/Ed75P6ULwaqClp2Ps7750JtynTorz/Pa3v03n8RyEDQHs+S6++OIk4Ilc9+Ljt/yMthP7Mh5B7B36/utf/zoJdW46PkSwezMB0P/ug5ByPukr7d9///2Urs4rzBBrPIHuWqz9OjjSUufAsxkGdx7vNae7a7hn7yhbqD0H8cqNyD3aLk29N37O3qH0IqLz7+22Grs/7yFmOPfgPef8G9Q6F+oh+TUIgs5CfcUtM0J2Bu2k7VE7iDiZNX80LARWxu8mDfIfzKJuu+22S0KNKNIo2/8Tn/hE+s12FsD6xpo1k08m8cRkz/rIosuaSXQTWH7Px7NaEqEEsHvKsLASX6736quvFosuumix7LLLpl4ZMc8qyrzvHK7FMk5ME339QUizmJqQqFF1HfdwzjnnpPufZ5550v1a496kB89LYK+44orJ6u55CTfbWX9N3pR2rN86H0SlSW+e0b16/vp0dtziiy+erjvnnHMmYel8zuve/OY4VluW7TfffHPc++CSwk/8jjvuSOd0XbhPabHSSislAQ2/5et6LpPO7GPCIz8jVm0Wy+9973vpPe2yyy4pHfbdd9/0LohgaeEZP/e5z6U0sW9+ftiPlU+HxnvI9/jEE0+kHqfr5/1dI6cHt4N2Ik35ufsENYyG+AQ1lC31hxGTIAg6C3UV7RHzF4J20lYhTWissMIK4wSZD+FTP7xO9BjCz1EPZGxuBDI26y0BPMMMM4x3DDG7+eabl99qgo1ll4g788wzk0WWAJtmmmmSpZMFfKGFFkr7athECiEUWYR33nnndE1Ca7bZZkv7TGjyo/3cD2HH+nvjjTeWvzSG2Z977LFHSgMuASy//idQPQMRzWp9zDHHpGdhRSY+iUFi2vHuky9XFtrEIqsv6+73v//9tJ2LBOHq+eG+nUca+F3asg5r4DfZZJP0O7cMEKkszCZE6rBILx0KnQjie6655kpi2zV0JJwvT0jI+xLC8Jt3pePCks1dw7vlVmNf+3lerhx8xe3fF4Tq+uuvP+696Ixxo+Gi881vfjOdy315PpZ12wlxfk0EurT9whe+kI5tN96J9AtqSOsJvcduRHroEMqjQRB0FspnGEOCdjMscaSJQW4Dma985Svpky2QjUCQc2/gNkBEE35wDh+iGRp5k8PQzPnhGiyhhG52V2gUFlKO7gouAckK6z6JYu4N0NjyZ2aV5TNOSOcOQH94lna5GLhXLhMZ92yWa7PphZz2JjpOP/3040LiSUu+adJSR4I4bvT89ut9j8Tst7/97ZbusVVci2tHDNv34D16N0EN6WGuA/ekIAg6C2240LXh2hG0kyEX0kSa+Hys0jnsir8Eb6Misl7gsniKmWzb7bffnmJMs8yyVOd9CVUW12yxnRDuIVtb8zX4cvNRZpk2aRLumSvIxFBgTZYzsQ+emwWce0S+RhasrPh8km3vL760e2T1dS5CHe6HlZqrQ7MQ86zXXFby8dmFZLnllkvfm4GAMJmTvzXrsGfSaTIZkP83ET333HOnyaUszq7FTzpbkKWbe6mHFdjEEPvlBVqIN9+5wgwV0p4lI4bte9ChkY+DGsqTMm5UKQiCzkJ9pa3JbXAQtINP/phD6wDhTkFw8pvlP0w48d8lRk2Cs/13v/tdsuaJ3CDChSF54oqLAmss9wERKliYhdLiz2wYn1XT+U2+4xKgoeKHy2fYcYb4CUDh6q6//vpiiy22SEP8BKxz8Ksl1Alu1mAT3NyP84hsYT/ijoATWYNQMtGNUOPfS9QRUCYhskq7jsKoIBKy7p/Q44pSP1xEIBL2jnU9xxHmzuMe690wuFywWPPtFrHDZDydBPfuPqWB+xQdw315Du4Tl1xySUpX5+ZKwfLuGNFApDV3DJMTHasHboEIaSvdNfQ6F1Zg0/BLI+4rJkpxsXEf3EA8v/TwDgxZu19ROViXnY/12fn18rmQ5Imf7oV1zrNLB9dxTzog0sl9Sk9WdZ0J1mX+457X757VpEfpyNXHiIO0cy2TKt2jCnHDDTdM98xVRIfJc3kekVac3z022kHrD+/FO3Rd+bXbUb69i3vvvXdcNJluR5qoS5TpWJAlCDoLRidlVHvUTHizkYx2U3vKjZR2Gikw6pl3R2MstdRS5dbBoS1CmngmoIgd4lNGdeP+Zt9WFlTfiRoikHAivgglgs+kQZmcWCbCiEd/iSjnf+utt5I4J5QIXj6//HOJWOdwbiLd+YlrQtfEQ9v5EhPp9jMBzXmILfdBhGVLMYHKb9l+BDAhqUEUes82FlTik9AzKdEQrnvwnVW3d8OpsLK+89nO59xggw2Sf3fGNm4txIiJibAvoenc7ovg59bgPoXj89c5PHt+RvvxEyYevQPPIV395j58zxZgx7rXfM+u792xIvtdGu+5557jrMm2sQh7ThZ/gpa7CsssCzqB7Z0Q0p7HuXSWHOf69lliiSWSX7b3ZjsrpvvwG8u3TpPthDTrP4u457TdvTu/e/C8+R7FnZZH+J7rNHnPzus96hjk79KxHYgGYiTFOY2CdDvegw6VjqgJw0GRKm2dLfkyJjQFQWdBXBGO2vRYkKVGCOmB07Y40kFrECOs8yy1YdXrbHToTFYl/o3AdDtGHLjacNMxIhLU8ohRH5OpGQuCIOgcGHKyYStGFWtEHOmBE86NwwQRIk4ydw7uE0Pp6xu0Bku0HjsLfFAbTTEqYhQhqCE9WLoijwRB56Gu4rY4kgRjMPyEkB4mDATwueVPKbxefxMhg+HHOxPD23sLaunBssN9J6ghPVhCIo8EQeehfLJK+wRBuwghPUzwLzbBkIt6vc900LkQjiZ7qoyDGkR0COkepAWfvMgjQdB5ZGOITxC0ixDSQdAg2bXD5M0gXDv6QnqYaBt5JAg6D3WVCfs+QdAuQkgHQYOERXp8pEf+BDWkhegukUeCoPNQPs1P8gmCdhFCOhgyDHtbqt2qh8IPDRb8U616KVRdO1EJG7aPlQ174OOvcxHU0EALixl5JAg6D/WVsLs+QdAuQkgHbSMLZdFILHxjkZQcIi3DUsc/bbCsmCpKi8DwP88rP7YLrgwRtWN8DJWGa0cP4puHa0cQdCZcr0Tt8AmCdhFCOmgbhrQtD27xHMHQLSJj6XMrG4KPsUVwrErZ31LorUKgs5AOlpWUmPYJakRafBz5PNIlCDqTqMODdhNCOmgLrNEEtADogp+zCG+77bZJXA8lLIJWrrQKYrsh0i1zzr0jqBGuHeNjBMZqqeHaEQSdh/rqvffeS58gaBchpIO2QEhb1Y2QuPPOO1OP31LlwvtZ5Q3cOqyAZxWlDKF9xhlnFEcdddS4z4knnli89tpraUWik08+OQmTSy65JC1ek/2eiTfnysfwu7bU6WDimSJqx/iEa8f4GDq2omHkkSDoPJTPiNoRtJsQ0kFb+OQnP1lMN910aU37Qw45JInea665JlmIrdpIaL/xxhvJWs1/GkT3bbfdVtx8883JgseizZL93HPPJcuv/w866KDihBNOSL7Xfj/mmGOK3/3ud0mA/+QnP0nb//znPxdXXnllcd5556XzDhaENNGoMg5q6cGNwSeooRx84QtfiM5FEHQg6qpPf/rTxWc+85lySxAMnGgBg7ZAVE011VTFoYceWqy//vpJ/Pqfdfn1119P+xDTxHPGpMOrr746LUjDqkw0zzDDDMXyyy9fzDLLLOMmJTr35ptvXuy9995JOP/mN79JgmWOOeYYt6jNCiusUDzwwAPlmQcH90+0D2bEkUkJ70aElPp32u3Isy+//HLqCAZB0Fmor955553i17/+dbklCAZOCOmgbRC3888/f4rasf/++ydBTFD7EBbTTz99scYaa5R71/b/+te/noQxsWwCom2iYrAYbL/99unvZpttVnzrW98ab4KiofMdd9yx+MpXvpIs0S+99FL5y+DC0ugegxoxsW58pIc8G1b6IOg81FVGSX2CoF1EbR+0BdbaX/3qV8VTTz2Vhs722muvJKh32mmnZHVmBeiNZdIJ64cffjhZpE877bQUOmzBBRcs95gwLH/8pvlb//73vx8Sq6hK2LP5BDWiYzE+0kNorcgjQdB5KJ9f+tKXBi1qVNCdhJAO2gIhbbIf3+jf/va3aZtev4mGBOgXv/jFtK0ex3zwwQfJcs3n2X777bdfMc0005R79A2XAn7S/KX/+te/Frvuumvxgx/8IE1mJNgHy/XCdWNBlvHRgYmoHT1IDx1K4R+DIOgsRO344x//GAuyBG3lE1VxEOv7BgOGmLr33nuLc845p5hvvvmSqPXhHz3bbLMV++6777goG3fccUeyVm+zzTbJx5nw/eY3v1meqUhD4/ys7fPTn/40hdHbYYcdigsvvLA49dRT03FrrbVW2r7KKqskkS6yh4Vfdt5552KyySZL9+GeTHysdycZCKKSuA+if4899ii3di/S1wiEkYHnn3++3NrdyCPXXXdd6kCK3hEEQeegrdEOaZuWWWaZcmt3c9NNN6X5TNpKbedIwbt+6KGHUnAAWmIwCSEdtAXWZRM4WJhVVIQt+DJbgCWHqyMy8vbdd9+9OP3005NVOeM8JoSsuuqq41ZENEy+zjrrFBdffPG474S2FQwtx8ySbbgu+2ELUffMM88kl4NZZ5017dsOWBn5Y993333FnHPOWW7tXrwrwlHHYrAjpkwqGLHQuZh99tmLySefvNwaBEEnkBcKU3cpo0GRXCuN7mrTRpLvuNEHHabvfe97xZprrlluHRxCSAfDgoqMtfqwww4rLr/88nJrbVb19ddfnyo5IriTcG9iZIvKYFJlt+Md/ulPf0qdmQMOOKDc2t3oWNxwww0pDKQJskEQdA6MNgw66i5lNChSuNmxY8eOSAs9X/iZZ545BTAYTEJIB8OCikykje222y5ZnzOsy6zV/J47DRMcb7311mQRX2mllcqtQwuLivjcOXwTC8ICCyxQLLHEEun7UKK3T0SrhIdTSMtL0uPSSy9NoxAELAuERX3mnnvucq+h4f333y8uu+yyYuWVV05x1YNJEyMLjzzySBpdyIgQJMzmtNNOW24JJjWEL3388cdT3aWMDgd51Er+qsdo6nrrrVd+GzoIaW6ZRoiD1vjkjwXhDYIhhmDmj/XVr341iSDDMD62r7baah258pQ+p8lk7ltkhuHA9Q3F8RfnS+6euJqIxW0hkKFGg0TIiv89HEgPjZL0yJNMiVmuPdyJhnr4VlrIx8R8rG446WL06emnny7GjBmTxJcyz23tlVdeSb7vI8mXtJtQPn3Mq5lyyinLrUOLvGVOCQOEPMUt0QRI/y+77LLlXkOH+kq4TkI+aI0Q0sGwkX2YDSnlD8tqpy7fSjRaXVFFXD85cihhgSbSTBA588wzi0UXXTRN9mOVtiT7UELEExlcXeaaa65y69DhPfDFt+jPd7/73bRgD4uh2OSs0zpkQ50m/MWlh8WJhqNjE7QHoTkNB4sCZHKzBaFmnHHGNC+D+47yFkx6ELGiSvnbX3SowULeUo+7B5Pmt9xyy2QIMdIxHAYaEUy0a+Ez3joR/i4IGoRwYzXQkA4XxPy7776bLPff+MY30v9mJft/qCGkubv0FSN8KBCG8J577klpIW45y47OGZcK3wmfoYYV3DuRLsGki3LG/98oR+4k6uAvtthixZNPPpm+B5MeyqfO/3DW4ZCv5C/C+bHHHkt1+HAJWfWoOitonRDSQdAgRBqrwXBOImPx5M/Gz+74449PoQTF0B4OCzkBa4h0nnnmKbcMLSYOcWux8mU9XF7M1CashxrWJuEe+4qbHkw6iABkMrQRjfwulX/vN7sQBZMeLMEs0cNZh6u7X3zxxTS6YTTxrrvuSkaJ4UJ0oYhCNTBCSAdBg2QfaZ/hgvWAW4eJMqzjfIGHM4IIKz1xPxwYGn3jjTc6KoJKttKzaAaTLqyW/KGXXHLJckvNH5/A5rYTTJp0Qh3OH1q9JZoE/2QdteF0A2OljxG0gRFCOggahGi0ouJ7771XbhlaiDPX57tpYRuL3BgSZNEYDjRKrCssd8OFe2AZ7xQ00Py2Y/XLSRflTBnnslRvqbNNWRuOCDlBeyBcvcfhqsPh2vy01d+iHVm8aTgxwkLYB60TQjoIGsTMZnEph8NlACy/TzzxRLHuuuumxl5Dn4X1cEDAGuoeDv9scOGYZZZZ0sTCDMuKNDJ5Zjj41Kc+lfwepUswaSLEpGXehbuTt5U1nUWrrIrEssgii5R7BpMa3HNYgIfL9Ur9RETLU9/5zndS9BftibUTGCWGA3naBO2gdSJqRxA0iMrPBJHhEI8q2Z/85CfFlVdeme5D7M/bb789iVmzvocj0glrMHFvqJKgHWqIVu9CmlitzHKwYsR6R0KUDcfKgtnixbfWCpvBpAV3KQtEETaiGfzmN78pHnjggTQhTKhO/vix9PukCzcGcyvUHUNdh6uXrOxrHQB5S5hOdZZ5HkLAGukYjg44dyVW6eGYnD1SCIt0EDQI147f//73qRIEIWn2t8qQgBpMXIuAFu6ONYXVTIO+zz77DJmI5bZAwFuEBe7Jffz85z9P38HiIvzbUMwCZ5Febrnlig033DA1Bj4aygUXXDD5Hw423gfrkjjW2ecyu3ZIF7gfIwcWHwo6H2VcvpZ/TKKVp7xL1kORYIRZDCYd1M+irOQoHepp9Xd27fC+fVevDbY7Vs5bYu5///vfH1dn6fD/8Ic/HBI/ac9odEUd7l5ARL/55pvp/6A1YmXDIGgQk9sshmLmt8gMjz76aPquMhTL2PaRjOc8//zzx03CEhnDM7OME7MmPnKrUCkT+MTHSEajbLlh/uqWG9bJEQ1ASD4NpfzCkklEzzvvvMUGG2xQHhkEwVBANJ522mlJrC6++OJJxOrY6uDqLBnBssKgekwc+pE+imTE5cYbb0xtl/QwUVtaqLs33njjcq+gWUJIB0GDqHAsO01IqngIJmGM5phjjrRgQ3/wZd50003Lb50Dgfyzn/2s/DZhWJsNQ958883JGm6SzEILLZQaIUOTwvJJF5ZijVJ/HQuW9Y022qj81lmI2mCp74mh6jT0f9xxxyVfR0JanGHhtfJIhQbLEK6lf4d6ufJugmvT2muvXX6bNGAVNcwfDB7mkFhB0MiREQYGAEaQ7B6nziK21eGbbLJJedSEEWbUQk+dhvpXvdwf6nCdh2uvvTZ1+vn7W1zIqOZwT3qclAkhHQQNwsJ45513pgqYFcPHUJkFG6yo1x8mlbDUqszM/ifCickdd9yx3KMHPtGWJ84xa4nwddZZJwk295BdBT796U+nxmEgsZyJPhb1/uC2kDsQJqiwZvDrc498pT2TSVrCg2mU+oumYTLXnnvumf53bs+kUevLcivNiFIWXnhu1ydcDb27NpcS59x2223TPgOB3/epp55afpsw9jv33HNT9BTD/u6HL61h3PyO3avGN3xrBw8+6TvssEPKR6+++mpxyy23pLIlf+aFLognk1Cvvvrq5ItKPHEN6gvlT35koXS8PH733Xen/GlpaWVxoEPxxI95D8HgwS8510vemxUE1dfqK6NJ6hP1h+gsE8oL9bBo/+hHP0pGFflMKFId5zXWWONj1mxugLfddts4NzeTkF2DgNUB5y+tntDBHmgkGO51F110UfltwhhFYwgiurUpru3DP3qXXXYp9wqaJYR0EDQIIZ1X0iOKNazEHVF59tlnp6geE8PvKluN+VVXXZUq+eeff7444YQT0tB/RoMvHBErsYrWdfndCpU000wzFaNHj04NvcrcOfgEb7fdduXRzeMaWbBPDJbrc845J02+IhhV/gQM1w4NifSwyABLG2He36IH0kM6Ej/8GE866aRxgqU3tl988cXJwiR93IuGSZo8/fTTaWED4oi/IyEuzvZAcA2TkiZGHhLdbbfdUnro0BBdnoXI13jLL8QXIR2uHYOHyWOELfFywQUXpBEFIwFGRQ477LCUV+QheVVHWF5R5iZkXfTODjnkkGLVVVdNlm7vmfVS/iKA5XeCaiDIP/JxMHgQu0aM5AP1FYODTrn6U4dX+WShFbWCi1Z/k/10mNXhfIwvvPDC1JHWUVYH15dv75ZgNeKgfnM9f+3DIk7IEvGu53h5aSDzOghk1+gPRhMdSR+uHazQBLV7bYcBomshpIMg6J9qRVh59tlnKy+99FL6Xq2QK1UhXalWqJVqRZa29Uc+R7XiqlSFWuXYY4+tVAVi+WsN56qKsEq10kvfq6KgUq3kK7/5zW/S8Y7F3//+98oVV1xRueOOO9L33lQFcqVauVaqlX36Xq3cK1UhUPnHP/6RvjfLRx99VKkKkcpdd92VzlsVm5WqaK7ccsst6Xfnr3YSKmPHjk1/G0U63nfffZWqYKlUK/Zy6/jYp9oopv/dR1Vsp3T74IMPKtWOSPrfPtJizTXXrFRFU9q3N9L23XffTf+7f2k8oX37w7lee+21SlXEp3eDqjCqVAVXSnPpXxVzKc3uvPPO9HswuEj3G264Ib2bRx55pFLtUKU8IW8+9dRTlXXWWSeV14mhvNmnKpYrY8aMSeWs2uGtVDu3qcyee+65KZ/6P+hsqh3vVB+9+OKLKQ94ly+//HL6DvXYQw89VKkKy/RbI6g/b7zxxkpVeKbyrbzvuuuuqW7NqKfVjdWOXfr+9ttvV84///z0Vz7cZZdd0v/vvPNO5cQTT0ztwFAgb6tr1dnuHdWOYdRPAySidgRBg1TLS7JqZUsla4JJZfye+7NGZ8QxNQkvR9rgTzzffPOl/zOsa6y5YlaDxZgLCf88FpF8LAsHSzUft77wO2stqznct4k3/ONGjRqVrBDNzNZ2r8suu2yxzDLLjItd7RqsdPBs0003XbLg9WeNrkc6mri4/vrrl1s+jn2yxYZFicXQBD/WetZ717MPi7176itqCCuz9DIaANbAquhKVinpwVWHX3OjeE+Gek20zEu0uwYrlfsycsHVxHBu/Qp5weBhUhkrs3djyF3Z8J5ZCH2MoHCNMmm2L2uwvMPayLLN/x9GnAz9c91h9WbVVCbVB/WwCJp8zMIJoyes47azjnPV4soh7+YyEwwuLM1rrbVWGilSP+WRplyHq8f4CVc736n+aASjHVwz1MPKtzxlxINrWUY9bRt3EnAl4UIy7bTTpuONavDrt498pZ6up9oRLF544YXk3w0jj0bqzNGRn8xVkbeMlPg0CncnczlWWmmldO9Qnzp/0DohpIOgQTScKkMVTz1EdKNC2n4aYz5tXBn40Gn0J4QKVcPee1liDbkKWaWaBXdviG+iOYsI17zjjjvSrG2N/HnnnZeGPpuh93O6P52LegjIiT3TQMniWQPmfjSQQtBlbJM+vfHuCGUiybvkgmJ4lvDhbqOhkl7N0Ds9XNc70WBnBjs9gr7J74AvtDxC+Bi+F52A4M0dzHqUKYKIL21fOKd3TJgRJfUQZzplXJ9ALJ1++ukpUkK9mw83sKEIDxnUyl59GVXu1d+963D7ySON4FidsByHmmhWvifUObK/fJWND/ZXb9bXvb07ZX4nri0CBHUVv39+++pu9bjY+TkCR6P09Zw6j7ljEbRGCOleyMD8O1V4nY7Cp/CecsopHxMzw4mCaZEMPoXDhcpL1IVjjz02WRvb0XCpkFk42rH4SRagKtiJiTfPodHvPaPa8QQ2i2hfaOzlDZPdWFxYRFS4/OJUyqzirMcDjYurcRjK2Lo6BKwn2dKjU8JCzufQuyZSCNneHQ9o/AjpFVdcMYlx1vgscHVGWIsmJKAaRSNpUiHrfTB8qIPkE1Y3ZcR7JnxZl/nKiqLy4IMPlnvXUEYIXnlhQuVKeTWq0WyEEOWYWCHq5Q+WyGDokQ/U30O5gJU8I2pIHlEzembCo8nM6qxbb721qTqUQUDeNvHccfXza1pBuVD3Ba3TFUKaqGD5k2n7+pjsZYJQRsZXEXcyWUQfffTRxaGHHjou4HyG0LJCl+fTMWANyfhN79Zvxx9//LhebztwbqLGBB8VxHDg3ZmpbciLaBRVoR1hpqQ5MUaoDQQWARNOWMdEtzCENyEIRxbU7M6RIQS5ZhCRfSENDAOqtDXaKl8TAU3C447CqqFcEH4DIQuWoYLY8VzcOkCw6mRwn5BO4lhL297LuLMk+t2HmGGtlz9WX331NGvd71wyCK2B4DzKonIQDB+swEYpDGH3xjsmQOT/erhf6NTquJrQa/icMSC7ash7DCxEcTNRFog3rj/KMEGl89eo9TNoL965+nsgdTgXEAaEbIGWLxhFJrSSqjaDpsjRY4ykWYBF3WwkzEhhMx14lnD7y+Ou26hLyoSQn50raJ2uENIaN76QhuxkaJESzMiWCTV6LHXZN5KwOPLII1Nj2+l4rr78/ED0qSyIA1Y6oq3eyk5IsFYSnBM6Ryu4roqFABwuiEZD9kLS6Wjsscce4/zBBoL01hASY+1AAzv99NOP86/tjevpCGh4e0OoeZ8TOlYaGP4jolleRSowlOj92GapY9vqO1jNkvPYUI7eyFs6HnyhMywzImesssoqKVpGX7G6pYdZ8u6ZZVAnxLObuS+v5mPkm4GgY6FxVL6C4UGdp74nOOT1HDIxo95XFnqLF4JEecp5RF7zITS8V4LH0LrjnCML7HpynWx/4kTZta8yYmSIfypf/Il1noPBw3tRpw6kDjdiwf9eHUJPMEoQ1TrwvVG32IfhI9fjNIZ5MbvuumuaG6KdEvWjL9Tz6hLn8de55F0ifN11103uQ8LoDQT5k6tc0Dqf/HGV8v8Ri14oi7MlXvUEiSpO/BpSFj0xFA3p5cklkwJ8nfSKDclo/LfffvvxfGVZPAz5qLhZ6VQeGniWFBYZQsTwFstdO+NHuq6hS2mrEWskNme70ZDpDJkExoXB5KB2dIxyJ0H+6ct1oBE0ykZHWMg18CpGE/icT4UsFqhKUqVrX8PP3jHBndFYq0BNeOGq0Rv5neC/9NJLx1nDNOoab/9fccUV6dwq6TzM2CrOoXHqqxFpFI0EoZFXTWTZ8b6IdILIvbtPz6UB1AHIlkYCWXqK50pAuQ/p2RvCSJmX3sq7d6mjQWwpH6yRWTwJbdYq3o178s5G+ippnYa0V8edfPLJya3LuyVarWQnPxkhu/7665OlWl4yOqMeJY6N0CkH6kv5R53hPapDjXjwnzenwCiG7WIQO7Y+36t3WLPtI5/qwGZjhlEb17eP+3StiCs+9Hjv6izuDK3W4YSw+iOvJ8DFLre16mQjsvZRj6lTdMDU57nzb5+LL744dcTsp43kZlePe8xzWuQf+Vpesk19qO2wXd1LBwi/2SpEPgYSfq/b6QohrcJjbTDzWgHgpK+iPfDAA9Nv/C0VML1MDeqZZ56ZKjkNoUpWPF+Nr4gHMnC2bubvrFp5WEfG5irCwq2gOE/vSSmo309hJHQN/REVZpWzmhu2NstbQ+88CqP7V4BMYnFt961x6C2kMypt+1lAwHAlEa3D4DhizHVVAuKr6tnqWfMPdE8El2t5dn6BY8aMSQLBeTybNGUNNGkuf1c5KZjiVBLphIuKReOi9w3Xdj4xiT1//s29EnvS23EmUoj/2bvCU8m4P+/Q8Ro1x0s7x+tYSEM+za6TrztQ3Lf0UvnxlW4F925kRB50Pg22iA7eq2f2rjWy8ozfWSG4Hog1msnbvZe+fP009ISB3x1LRMg/OjYstvKr9ywfm63eV/5sBPfsWjoAvV1PmsHzyGfyo+FPDYM8Sex7n/KshsZ+0k/aGx6FvCY9Ha9T3JeIto/RFyJGg6NByx1JeZ1Il3c8C6t270atGZRrnRgiLoT00JLzkc6Y9+u9q5NYgtXxthMx8hc/efWK9+59ESrKiv0zjALaBOWEWGK5k/ecV11MiGcrI5RfdZl3r2xwHyG03Rex5HxGQHXuWSHrrxUMDeoP70m77z21ijykvdVZ0ibyufc+vV8WY3lLnnM9qItzfUAIm0joeL72fdU36j551b06jr6Qj+Uhrnnqcr9pYxkV8pyRVpCv6R73GLRG1y3IolLj98Y3svfwq0y/7777FmeddVZyeVDQ9ttvvyRU+SHLuKwZCsmss86avisQBLoJfxpR1hAZkyj0GxHTe4U0vxGAllHm60lA8Pt0HRW2e9D75D/LkmEWOOsqyzEBRLj6XSFyzwQpwaGC7g0L20EHHZQstAcffHCaBEhosmS6B8cR4YQvX2rn4Fvt+flPa0SIdgtf2O4epKGesaxDlKsYfCf2iG+9cMJdZcCaIz30rD2vZ/KMQpBJP/u41uGHH57SdP/990/7up4GS4NXP1Kg4WMJMIGQddXx9rcgieeQ5hbn4Bdt6EvloMPUDlyL9dNzuq9OxfvQSZOP+upctQv52LuUp7y3TkU+Y43WoRqI9b0RNEjKicZtIII8mPQgqtQ76sjc0Qs6C3UBo482rC//+U5Bh5BOYQxqdmJrszDauRb3uKA1ImpHHYQhq1UmW6nAKsbf1rAv4eA7v+Mf/OAHaZhewWT1IrgJXAJG79FwNYtHb1yLn/YxxxyThB4fJYKaWCMgiRSVMQHMHYOYto0llk+3a5vQVz/kPzGIPz5ZhIRjCd8MC6uOBWsluAOwkuaJbK6r0+GepYnjrdDE6ks45O8EMdEM++r1b7HFFuN+9ywqCMPwxK508tEBkQ46BYQ/K7R09Xy93W38Lk0JfMc4N2uAfbP1WXp6P5YMbpeIhkqNJWBCk0o6Bc+ukRhMEQ3vN1uLOxmWIvl+KCwuyhILt3QJugt1mfqq3koddBbZ5aLT63DttbY9u4MMJvJrX0a4oHFCSNehkOVeGdFEILCs1m9XWebvhIRhcRZAQpobiN+JSYLchILdd989CdF6CGxCldghilmD83aimRg0VC7eqWtkQURo8tUzfM2lguBtdLav87CksxyyGLM2s2r3h+MMZ1rClKvJzjvvnNLGcyvs9d+lgR4/pJEJFIZGCWMWXKKbhd1QPKEhnXQa+K0T8obZuRp4rgn53Nqfr2GO2uAeLOThfCwNg4m0MKTX6SJJmvTlOz0YeM+DLdgHinyrTA1FSDplWFmQh4PugqsQQ0urrlLB4KOtUn93eh1O3NIP7Zjb0x/a58izAyOEdJvRWLOUZmspl4zejWq2XnOl4F6RxWd/OM5QusqgFTTyrM46AXxoDXcPBazTLNqEqI6G+2AhzOnEmmyiRiNkq3i28ksL1mliTvoMJjpEfJv5rgW1d6FTxtUmqGFEiS9u/chWEASdAUOM+jvq8B4YuOiRoHVCSLcJgs7QMR/mHLOY4OMv6W89LMtcG0S2MIGAkAQhOLFQYgSoa/Bnsp/9uYRwjeD3nN0qJgYLIgswa3deKhlErkkN+RzuUcQI528lvI57630uE70MqbH082U2MQfEh3RqBL1ny/6aiGiRFeLWX9uza8pgIY1YClilm4GoOu6445IffV71DPKFiZJ+40fv/3ZD6PKpN+Gz3UgP+cnkxVZwbyKL+JsxWUd66GQ2mieaQYdO3jGJdzDErjJqtEi6BEOHfGOSsvfK2JBRt/ABrR+tMoJoX3NhjI61G3US1zmTsk0eDjoH5VM710wdLg+ZG6Ve4gNvPlNGG2fejMAD9XV7OyH6zYMarHUZjGAyRgWt0xVROzIqOP7NfHSJONZjDR5fZNY1bgcm1nG34FepwIkMwcJkKMjwh/Xt83eiKn/3P/cEoZaEttFIi5bBGi0SQD3uwwS5LCD4PRNRthOujhMdwlBhbiD4T3PN4IPHvYMV0ExzFbZGwhAQt5A8fJ2t1wogEcvqTfD4uCfREYRock7D3kSR6xPkhK97ItbdI79gaeKanluhs4hLjixS/10FJRKF60tjlYBjXWvbbbdN/qOEhgbGAiGey3456oPzqKikp/vqjYqQ9VmYKbOjudM4niuDmfAmTwohp1Lzbr3Tdk4wI35Z1RutePh0c93xvNJXB0KYIcf7TV70rp3X7O8JxYVuFfmQT7m04jbTbrxnZcd7bQadP3nMPIG11lorpakGS5hK4sb/8prhzXbiuvKO2Oo6lK7bTvKICXeooXAlCYpUtxCtypb3ydiQO3dGrogc9ahRLx0po4CMGP43wqQ8Nts5nhjKhPPqJMoLjCVBZ6B8ej/a9kbrcG26hXq0JdpE7ZOoQoxn2m0hOtWz8qHoGe32v9Y+MCqow80dajfaJe1qu9uebqKrhLRCRNAQMASpxpp4yfE8+Qz7nd+xXpqMRYDa15AQx3+hvuq/s4b6TnzyXeYXzOLh3CpRvsW9G2sFUGEz8S7vJ7oFMctaa3/nVtgJShMefScgiUWixbGuyTrLt1h0EQI141nt43n4KRMQxCpRnK3Pwj05v/O5J8+rwXFPjnfvRCj/ZgJf2B0FTlgnApjQ7f2dSJd+7ksa5RX0iDjbsyuGe1YxuZZtJgbmwPbS0DF9rR7meiZGuFeNpGvoCO24447pGMKdEHMvrNQ6RBMKdt8s0ltnwftodHKG/HPEEUcka7R3R/ib3e/+dEw0tjpg22yzzaBUZNLLu5Ym7RbS8oj3RZh4382g4TEqo1HaaKONUp53LqMzxLMILI36/zeDPCH/Cfc4GEJaHUKo66C2+9zBx1FfcVEjopUheSmLaEJZZ00dKAITIZ0NHSL6CF+n460OamcMXfWZ9kPd5BNCunNQd2vL1Mva/kaQj9Sj8pf20iR77bR3zKil3hY1iouEvNaom2Kj6JATuwxngyGkszFL5yBoja4LfxcEraJRVHGqQHV8+oOwV2kLX8QHjRAnOoVI5FZjCWKVsg7P8ssvn0RAb1T8wiKq7Ahi1luuPTodOlc6b+7JgkKil/jrnO5RR0TnSTQVYQnHjBmTRIPvhDWhpwEgao28EJlCOeoYNTL5xPO5HouMiDCN4pmMkhA1RiB0JnSGnOuMM85IHSzPtvnmm38sXrcOIfHjmVmsde50DH3X0TQ5mAXHM2rQiGbWHKMT0sIEX9FdRJMhqFiQdI5YKD2zzoZ0MSrEAiQNNWLSpRF0orlCiXiTO+jB4OC9EADCPOrwEzc6dPKE37xneVP+UPYsyGX07thjj02jfDr93ru80jtEqU6dMqps6BTpBPsuz2fjRXaX0hHO7nYMJKuttloSXkaiDP0L+ylP+u4+jB6qP5RhI6QMHcRYuzr8wYTxPuQZ+aOvmPP9oT5XX+nsyxcW6VGHqh/U7VyLjHbVj3AQ2Op6BhTHyD/qX/WdDpyOlg6fes8kevlCflIfMbjYhzuaUWyjizoBRnnVg4xg8p+RY7+Tc87HqNaoZZxxR+ffiHHQGuEjHQQNwtKkImwm+L2GlwBXAcM5bCPsVJKs1RZrIL5UtPUQjQQdNxUjHxpyvnqGELngEIAaZu49eRIkVyPCnIuEfeqxb640nYNvnwqeCxBB4TeWcxV1o2gwmgkrZ/RFA0Lk1K96qQFQ+Zt8KhKM9NJ41CPdPCPXHc8obfyvEdHw6AzYh/hhoSRedB7y9XRg/JaxLzGfFyIisrLPtnkOOi86IKxMjaIzQtC101Ug6Bsji6x0ypTOj9ENLh7eJcFEaBDYrIiQ92wnoIkUYtfHe67HPsqDESNlUp7IbnSEkv2NPDi/PEaY6cjJm/xYiaJ6lCflzPHOx4Kuk6ZzLc/pVBJkweCj3lV/9+6gN4o8pIxb84BBgEiuXxRLHZtdNsGarc7mxqielT/UW/7XsZJ3tA/ylDpKvaeDLw/LFzp89TCEcCX1m/wm3/nIn/IYVxNtgOMbRdlpNIxu0DchpIOgQQgvFRTLQSNk4c3aLIa2RVJYR/mn+40F1bCdkFnCIdZPiIJKmNWLlZTAFEqRlYE1leVVhU4IEG577rlnEscqehY3C9qo7OshPFTkLGdEK6HOh15j4NlYVVhtG7FGZzQm9ZO7+kNDQER43no8h/TQ0LkPrh2sLvVocBxLdEsPoRwJJRaYPfbYIw3pS1d/N91002TlI6jFf+fBxgLlOTPOp+FhwWe5lnbEuPTgNpRXPmzGx15DqlGULsHgIj/L896/YXfuXUYEdCK9P1bHVoarnZOQZkmWd7i4KXcWWmExlEeN+LiuqEzEkDka9pVv613soBOs3LOMczVjjSR+XEe+Y6HmZhcMPsq4+ltHvFnUXVyJ5AV1biO4jvet7pE/1N0MD9ZVUK/LS/KFelc+yx19dbg6TVtRj+sT0cS0+lIe0ulX36jP5CUjHNm9qRFck7EhaJ0Q0kHQIAQccduMSOKOoXHlo2nIzvBbXugmozIleutFHlT6BIGKkeA2hGfYmrXTBFaWasJBQ83qptJmWWBxc77eQ3XOxwJLbHoGjbdIKvy9HedaKme/N4L0cE6VeyN4PmnAN9qQu6gJ7ofVRYOQkR6eOVsSM67leTVi9tHIbL311kmc+J9lhfhmWbcPy6L9PJPGjwuAfTLOx6KoQ6IxIbx1UKSvzg9BzZro/I3iGVmknDsYfORVFkYdVu/WsHm21LEMm2jIH54V0KiFPOXdeN86Pf46th6CRL5QZnWmuEzpULFicsngauU479q+8qS8owOqbPee20GA6VzpuCqb3ESIKUP28iZh10znNWgd70zdpxPWLOooox65/lYn6zR5//KUUQrvV52fcS31kLyk00RQm/thrhKDAUuy0UT5TR5wDnlJvSUKFeFdj/uWX4hv11TvyW/cyNTj7jGPtjSKfOkeg9YJIR0EDaJyUlkReY3iGIvLWJ5dw0kM9/aFVJEZ5u0doUKlrCHPYfHs53/b3YcKk4WZaHQd37ltQAPfO76zfVTSrB8sHu7J/1DBE+mss4agG0Fl7prNWNPcO1FCfKu8NQa9hSfh4R56hzN0LJFLFMF+3FvgPogcs+s1Xt6RfTU6GhfnJ9rrBbvzadA0clbAZLXmbkKcafRYIFmTCKdGIbp1Ynp3AoL24/0qB/IDYSvP6/gQqTpOrMbymc4vAaL8EMOEs/Jm3+wHX4+OlfyUY+sSN/IBn3zzB3RcddhY/+xLUOV8mPetR55Q9lkglbuddtopbcsdYnlQXP9mhuOD1vC+1A3N1OFQd6gbc4fNSFcesTICIi/Zx9yO+rIvDxLFOU+o84wI2kb8Ooe8lPOr+5Mn5Vl5ibuH/zP2ySJcXuL3r31RtxvlMwKjDXCORmG9lpeD1umqqB1BMBDyBCZWDYK0EVSGJjLxs1Uhit+tEvc/H2ZDyCplVgzRUerJlmEWXBYtFXYeBvSXcCAc+RRr5O3PFYTVl7hg7VBZm/yi8taYm5zCb5j12j2xhDgXP1D3StQSpCr4/mCRzmKkEfcH12HBIdp9VN6eX4PgehoA/qNcXJxXehA0mZweRAfruQZIuoiaoyHxO79DEwp1LnxnQXJeosiH8GKh9JHmOg/STFrppDifiY+jRo1KFmloGA3jNwLBJj00uCGmBxdixMdQN39lYsV3k3t1VuUx8xBAQG+55Zbpd+VXPuGS5H8Ct/5dyUvKAv945d0Ih3yoLMnzyo78YnKwzpiOmxEW5+PmoYPH2m2khTjOgtt3Ysu9KruG0/nO6gQoGybHRp4ZXKS7+lGnqpE6XAdceTa/wjsmeNU7OuhG87xrdYn6VZ4RVaN+Do38oS7LdYwOl3pJZ09nSv4wsqhdMDrhfNl1Q17yu46aOjuHalRvOZ86UB2us+h5tBPaFXlJnmu0jZKf5d0JrSYc9E8I6RGCBkFBU+AILT3XVtBQKLxmBxNdw12xE68EkIZvuGe1q6yIWZWdCq0RckWrcSZ4syVEha4RVQn6bfPNN//YO1MJE2QqTPuBBYtFxDEqVGnDHUHl6V2pxFXC0o1FV8WvIWA5UbESnd6xxkSFLgQYi4T9vXdigbBoBHmOhdcwem93lUZwH+6bJd7zsEK7V9v4nPb28Xa/npHoth8M5XNL8RuUgSzAiRfPTEx7d9KScCa4/M8iaJidhSf7eTuf4VKCy7mcR3pIx0YginQO3FMzfopBa+hAKlPErrzBDUNHKCOPyRvKhU4U8WK0wfu2XXnqPVmWcJEniCMdI/lE58yxOZ8RWES6fKJzSEQpC8qwTpffdVKVJ/lYR5Nwdj55ysiU8q0ekGfE3m+0sxa0jvekfmQwyKNxE0O9qK40CVDn3PuT59Sjvstz6nhiWfvU+x3KM+pr7zi7b+gwyTN+Uy/pXOU6V53uN6JbnUjcyru+y6fqM9eR77gw5fPJr87lPoyaqI+dvxF0Fhkv1LlBawx6+Lv63r9KyDCaxirj8jJEXsVM5ll11VXTEElfOJ9eGP83zviZvL336kIynElasI/hmTwMV/9bRsERDsk+7sX99rVinnPlGdf2M6RCZGWcm3+TQsfyKIPn7Sp7DXkzuC/XE2IHzkMwZAHlHg466KAUTsm9azRaQUVhEpd7JgAJj0ZggZFueThUIVY56O0ScQp8s0hjFZiJc55bRTScqKhYj6X9YK+i2B/Sm0A0zMyfdzjwfogH70Zc3uGGr6KJN1tttVW5ZejRQOsgqeNajQwQdC7qcXUAI4N6LZi0YLFVb9Idw12HE+CMB6zbRgGHC0LaKIlJ70FrDKqPtMxKXOkByiyGToX7kpEz9hGGyzCqj/300vtCw23o16INfBrr8ZsGLJ+HgCNy7Z8hRvk75n18+kLvUWVpcpLoAH1ByBiy52fqPAoooWfWPzFrm3vyfJ7JCnaWPbbdsc1AwAm75F7yfbuWoSbD4ixsLCDtmDDgfrPobxTiW0SKM888c9z9EXiGMt2fHncruBfPzorQCei06LCwJA0X8o4hP3mPgB1uK73OMcvvcMJaf/zxx6f8xndwOJFHdLT8DUYO6iBtmSg3LJQhoidd1N/q8eGCgGZ0s4oyo9dwu1RIi+Guwyd1Bl1Ia/Q322yztE49LxKimo9jhmjjl+h3H2JxQo2h87H49FUIiF/DLfk8Qs2YBCUMFoha4rh+HyHJeuPcVjwTTsy+JnOJA1mPc+kMGAqXAV2LFd1fxxhqcW5DNH43IcAQsklNthvuaxTin4+nDojh4nzvvluZSZqo2LMP4EAxNGmSVaMQdt7nUUcdlSZq5fvzrj0/QUFUt4J3ocGyCEknkIf56iesDQcqYuXA0CK/uuFC3iMwspvFcOG96LzpgHeC+49hWB3rYOSgzvdOGSzCl3TSRXul/h7OOly9yfjEt55LRr1P9XBAgzU6wTzom0F17XDqHBQfKiFO9Xx4CEqVE5cOE53E5zQkWx+eqi80mvYXN1RmhOuwSvF9y99ZpAkwVirCVQNHIBPphnT8PyEcz6XAAhg+BCv3lIzCaDISkUgwEvHQkHMV4dZgYYuMa7PYjh07NvVAPUO9m0aG6N58883HSwOFzb0ScCzuxGlG+vHj9BsXDBYTbiPZtaP3dXqLZPdrQQsFiRWNjxRfPdEevA+uHb5bfY5g8t7qlyiVTqzNhvWdW3iperxv1nLppRPDYi5t+PTyHzVRjmWdn640NkGOy072adxkk02SaOT3zfKfXTukJ79cbiTum1sNFxzX8bw6PtLD8/WekT8QXNe5vafhHhbsBOQ/DZKRH/kuqLl2WBiBoA/XjiDoLLRjfN/VXfUupt0M1w6aodG5McHHGVSLNKHZeza/Xn29TyexYzIG32aWTAKpWVwni2gQeKxk/HLzTGsNHEsCsWUVKbNwTeKaGESaWLx5EQs4l+OIz74s5woosWWoOX9OOumk8UQzgUt8sKIR/PbnqmI2sOMzrmUfApWwrRfRIDhZJVnAe+MahKZYvdnVwv/iqkK6WwGJeGVZdw1ivx73opDpNHBPyR2GjN/5vuss1QvsjCE071+6E1yGRYl9Atv9EdmuL08Q0DpV7tUIBfcdnZneELPOYaRD2plkZBRDj5rQNtPetfjCS/t2Ip+ZeMTvPaihjAynVbzTMIqiIzyc7j9BEPSN8qn+jjq8B4ah/gyYwcQZVCFdD1FIjLLS5NmhhCABRkAfeuihSawRUP0J3P4g0ogt7hYZ13IdPruc6vksE3YTQ6FbbbXVktDno4x87vrljevxnKyoBGH9h2U547xm97ofLho6AWbZmixYL5adi6U9C+ZmIDjPPffc1JlwHWJTuCaWXW4pBLCwaCZs+j3HOc5kIS6dtttuu3S80YR63J8evvubmLuKWfBWCbOaEyFKeOVn0oHwV+eGFT3fqxXDPENviG4uNISzSAoqRK4vrOc6BHzPLIBiRn2jEyUbRZoYATA5Nqi9fx3U3vGquxlln/ta705nEATDDwOS+jvq8B7oEwapoHWGTEgThCYVCgFWDxHJ0md4nqjkrjHQl+pahle5DKDeYk3EciHZb7/9kkV2YjiOD5PV08aOHZs6As6tEPZlBYbz+40gzB/Cr94Kn/dhmeU6whpPRPcOiu76eopZsDQDEWoyYp4NzKWCkCZkWcdZg1nNhPpyP4a56iMhqnBE7nB/E/OZdj73159wcH3xXV2X2PXsRg1c3yiBexKXE855+OGH9+mLmN1EWMNFaSCkd91113H+wsIHmdRJzAht1W5YYH2CWv7UIfJugxrShIVHugRB0Fkon+rvGDHqQfuvzgpaZ0hqe6KHdZSP7cRm1fObZUmsd29oFscKgyfe4oSspBo5oo2FsT9kMlZplvQzzjgjuWG0w7fKtVlSuR8Q9X0Jc4We1ZVFnH9076gcBKzeZG/f5Ayxyn8azqUz4SONXH9iUT6kEQux55/Qym5+EwbKJMr6CaQZ1+GmwQ3Dvt6/RRJY97mM5PitnsP9sG43An/sH/3oR+M6KoccckgS0N75PvvskyoFsXz91pd7SKt4BmELh3tySCeh0zOhUJXdiLxnUrB0CYKgsyCi1d8xf6EHxjptc9A6gy6kiSk+woQZNw6iiUWyL1FI9BF8jQRKnxAEGesx14AJ4Z4IU64G/eF+LADhfM5rMpu18geC67O680kmykUWIXr7EsSsfdwvWGxNYMzpJr34CLOq9yVA9bi5NrBKS1fX5CdNDOqscOMwDM1yD+nG4p6FN7G6ww47FDvuuGOyDhPDvZE2KiSTAm+88cZi9OjR5S+1Z+QGYZJmnhTqWbjVsMBffPHF46z0xIfJe6zfGRZ176g3nkuhF2KQlV66sT4LrchvnSWdgBYphYsQC3i78EzcR7ggBTW827yYSVAbMTFilfN8EASdg/ZC/R11eA/0A4NX0DqDtrIhoSeiA+ujBTVYIk0o8yEK+UkTUER23k4QEZYEoOM1SHxn7ccSSMiYREZwEaKskCyiebEPx8gQVuUTA5pvbt7u3CJUuI5JfSamCRfXe6IUQekaFnYg+O1HOPNdFmWCb7QQdwQi/2ECk/WJKHVfxJ9jCF4dAsLV/TgnK6wOhfvm7mGZT+ci9qTJmDFjxoXry9if5ZZo5JtNDLum5yAepQ0hS7Ty+bbN+a0Wx1LsvARydqngm03M6oXmCYcqFWni/qSHpUZNApSu3GNMNiSW7Nc7vBhhK0Qd4WCyoL85jV2Xa0z2VfcsLOLuX4UmLGLeblEZHRWuM45n+c/p6r3x63bP8obtorFw7eCfSzAvueSSqULg1qEzYBUx98a9wz20A/cstJn7bdZnfSSiXOm8KFvt9kefVJH/lTVRaGISZhB0FtoT7YN2PurwGvSK9j0iUbXOoC4RTniJTkEsmmyXP/xiiVMNMYtp3m6p13orMbcFx3MxyNE3RIjgj+ucGi3h2eobLOKKO4TfM44j6rl8uA4BKdRLX0PS9hUKhjhzHgXPREBCmrBkRfWX0HQuAsJ9GC4iHAl7LgaO8xuhy+rrGG4ttruu+/G7oSbnsd1z9rXCEUFoO9cXx9nfNT33brvtlu5ZWhObrM2EnvQl5N2LzkW+R/vncxLFXB9ymoiwwVJNcDuPjohY3K5DvLISix5SD6u0Z3N/rNj5/pyPmOg9QVFnSFQN58mLGuhseL9E9ptvvpmO90w6Os5nfx0sQta70LFwb56ZBdA96iA4Jr9r2z1fK0tXTwjn9p4I+naJ80kZ6eGdyBexQEUNDbQ8otxFZIAg6Cy0P+os7VnU4TW01ery6Fi0zqAvER4E9bAacxWxDHnvcH6djgrHiAMXlXbGp55U0SgZNTKywg0oqE10NlJlhIRhoJvg9mT0SAeCdUtnPOM37l/mm/QWMDofRtSMAmayy5jOspG+PJlZZ7uvcwRBI+QoQ+ouZTQo0qR/I8hbbLFFuSVolphaHgw6LAAmVvIJ5+rDMj+piWjocwq/x2Ie1NKD5Z94DGpooLm7SJdugtDlRmbeBtcW8yWy+CWihbQ0dyHPwaiHBd9onmN9hLY0ByL7mxPZtvtrnYG+zhEEjaB8qr/V40ENBiJ1VtA6IaSDQScLUI2hxrW3u8ekAhcU7jf1lkbPpmLuNuGE7NbDtSaoYbRC2EY+/92E/M9dTBQiE5RZkomW/Js5IxNKE65oJhDnBayMVklDZYs7m++2iznPxWtC1miWbYIgT77mckTEB0GGqyW3Ky6Y3QijlrZY2cooY71D7wbNEUI6GHT4gfMt1xgOokv+oKPy0Ujnikijfccdd6Ql1Osrpm6CSDIvIaiRxVy3dazMG+DuxLps+DxPaMbUU0+douhMaPKl+Q45FKZ0U8Z8J3oInnweIoD1zMTzvpDuFmYyJ8S+5n9wNTF5WvhVlu4Q1t1Nt1uklS2T+blLmZCv3VKmYlRxYISPdBA0CJEgXrbGXuNuIiyfaUUor3zZTWiUwkd6fDRIfIFNpu0GH2kTjHMMWqNNyoePScssyRmRXSzGJUrTxEYwWLIdzyIt8lBG2ePbyp9z8803L7f2IC+aiG7lWh8jJdxDTPTWkedbbQRFpCCTvUXfCbqP7COtw9t74nw3oH6yLoR5HCbi8xPXYTXJf8899yz3CpolhHQQNAgBLbygWOJCIRLSGmercg7GKoqTAiwcxPRAYr+PJLgTsIgKPSkywEjHpEArv4JFWCdCqE/hKwlirlBoVEjLS6zI9s2WaAjRdd1116WGv69oS6yMRodEgRLSkzAwAuZawoZaw4A12uquEJI06D7U4aKBoRsXZfH8OpzENAFtsTdtl06rSGZBa4SQDoIGUQkJDciiQSyZXCWeuXCOvZe+7wZUHdw6XnzxxZgBX0LQCZ9J7LGCjnS4a6ywwgrltxpcKqzWus0224z7rREhzUpIABPEvcuT8nbppZem8/aF+PoXXnhhcgVZf/31UxQCC1hZw0DMeX6gfGOJBr7cxH7QfRjZkJfUXX11yEY6wuAaRbXmA/cpKyr7KzSuchO0RgjpIGgQlfBtt92WhrMtKMTXzGqUKicRCQwhdxOEj0D+htDrh/G7GdYujdRKK63UtXFZxXE/++yzk4Uru2c0IqQNu1v11KRe6ZfRgdVh1XHtq8PKrUPnRR4k3rmaEMrWDTCxmb+0Tg2h7bvFwYLuxKiJEUV5pj6PdQtcO7jiabus/WD9BSM12rG8xkTQPDHZMAgahBuH4Wb+l2LlapBFElh33XW7crKh9BClohuHSCcEa+cUU0yR0qWb0BhbVdSH5ZhrS/ad1rkwuYklkOuHfbM4NlE3R9nwlzXbwlD12M5SPaHIAjq4OnT+8n12fv7ahq4J7MsuuyxZ4ZTbbuvsBuOjkyYf+HQj6iWL1R188MHF2muvncqpyb4s0kHrhJAOggYhHPm95qXnQVDnFSy7EcJkQtEYuhGh3DTSBHU3werLj9lHp7I+aoffpIttyonv9uEGY3KhkQ0oS0R076gc0pLLhlVse8OyaOVTcah32WWXZO0muC3a8sMf/jC5liy22GJJWPPXnph/djDykQ/V3/V1eDehjE0//fRJQGeUyW7tWLSLcO0IggZh8RJei2tHb7/QboQAskgGa+O+++5bbu1uWF/Hjh1brLjiimmJ/GBwMbnTnAVD1TE0HfQH1w7zXNRdymhQpMmHotvoiAatERbpIGgQFunPf/7zXRGNoRGkRw4tFtQwdMxCHy4EQ4M8yLVo5ZVXLrcEwYRRPlllfYIaLNIxqjgwQkgHQYOohM38rx8W62ZyxyJC3/XAB5FvsHQJBh8dFm4feUGXIJgY8ouO14QW9elGJptssq6MYNJOQkgHQYMYDrQalKgEQS38Hd9T4e+CGtx/XnvttZQuIxnPZ+KgyYWiYeTnzZMIbb/44ovTtkyekCjOs//bjbQXkeG8885LLkdB0BuuQL/97W+jDq9DCNOXX365/Ba0QgjpIGgQwtFEKZ+ghslelpgNasgjGmvpMlIhljW8BLSOpQVPxH6GyYZW+bSwCr/lu+++O23Pi7XodOVj2400F0/66quvTsuBB0Fvog7/OAxE6qygdUJIB0GDcO0wJBjh3nrgLx7Dgj3wNzQrfiT70YubTqgK83fMMccUq666alp1kEWYNfqPf/xjccIJJxQbbLBBijH+l7/8JYWlE9v56KOPLrbddtu0X7utxvxerTI655xzlluCYHyya0fU4T2IrpNDVQatEUI6CBqENcOiESN92L4ZWDIIp6AG646QbiPZwiOEGEEivrN3zx9caDllg8V5ueWWSx0KvstC17FAE80mNE099dRpcqqQkZbYr0faEdwWbRk9enRa/Ijg9p0Fm7XZ72eddVZabEU6n3POOen3Sy65pDxLD84n/rTf7WdRmOz+YYlw9yqCQ9A9GLVQf0cd3oMykZdND1ojhHQQNAgh/fe//z1Z5IIahvkN2wc1NNQEpXQZqQj/OPPMM6dycPrppxe/+93v0oqBXHwIaxNykSMkWIjFimrf/va3x203KbO3nyphbDEX1m4LqYwaNSrtwz3k3HPPHZfXCGHXvOeee9L/BPJFF130MQu3exGKkAB3PqstckW54YYbksD214puQfegcyXfimEe1NDpN2oUtE4I6SBoEJa4ySefPFU8RINKudvhwsCVIajBUss6O5LDa7Eysyxb3IQwJUYHupKjssSvmvX6+OOPLw499NBimWWWSa4ae+65ZzHNNNOktOVOsuGGGxazzTZb8s3eZ599imOPPbbYbLPNxvPVdz6rJFrVUJQdx9qf6CasDe0T/AsssEB5RNANyAfqcPmo28n+4jrGEYlqYISQDoIGyUL67bffLp599tkkIkyyeuaZZ1IUAsPQrG+GylglR7rVI6/0OMMMM5RbAi4NFmIZyT7SBCuLrs7C3nvvnZ5VpAzPLpSWCYfIbj9Eq5XTWJHzdhbq+mWJNejKDEHOZ5PI3WuvvYqvfe1ryQefD6eyRhyzbCtjVjQk6ImijTbaaDxffedjvbYf4Uz8b7LJJkkwLLHEEmkb15QIU9hdENLyVLcsiW2ETDukLHDfEFGIe5Q2THl66KGHUtSOMAoNjBDSQdAghDT/ThZYFY8PQcCSZmjMMsWPPvpoEgzE9a233pqGqV999dVUYRHbRAaxPRIs2oQ04RPWjB4INsKOqBypEKBPPfVUEqssxpbivvnmm5NYnn322ZOFmhuGcmAY3ZLdrPTyvjKgUX/66aeLRRZZpDxjzd2DZYzwto/jhSnzvzL3ve99L62gqbwRzPLdF77whXGhF7lcsTZnnI+oJ8B33nnnNMmR2HYNE4a33HLLdH6uJEH3IF/Ip3n5+kkdVmVlRSdUfla2iGTtkHbHHACrFmbxzNijHBLPOpPKp+XSY/LlwPjkj6uU/wdBMBEIRw0xIW0i1Ve/+tVi1llnTVZqE6myFdJ2VgCVlW3+Z8HzPyFgSWNCmmVOJacyU8Hz8SSu/W+b/1lQOhmdi4EO648k5BEiWrqMVFi5iGS+yzqRxCzXi9VXXz3lV5YuDbd8bhnm+eabL23X0HOv8BtL8HrrrVeesZaPQAw/9thj6Zw6phb7IaRd85ZbbimWXHLJVP7sTzzzgVZusqB2PyKIKDuid/ziF78oHnjggXEdWqLhiiuuSNY5IsR5TY4MugPlU2fXZ1JBHtVp1WYQwT7aFKJYfteOcIkyn0D+Vs6UT2XMfo5j7PCbtkmnlnDWdnGRYqHP8xqC1gghHQQDILs3EJMqKcPOrB2EhUqKyDaMyApmP5UZC0K2wBEOGnSVnoZeA28fQ3AqSlY3IoAgsD9rIDHuf9ceyYIt6Ex0FDTMrGAabEL3Rz/6Ucrr8qWG+YUXXkh5fosttkjHKB+2E9csgltttVX6W498r6woE1wyNO6LL754+o1YkPdZpl3Hvs5nX9tdd9lll01WNuXLPvPPP39yO9KJJSZ0fu1DZLN8Kz9rrLFGrHIXDCvqf/kzuwNqA4xaytfKF6uyTiNrszZB2VDv60DKw9ob25RD5ZJRx0gMF7PpppsurfqpPGifjJYpO8rwSB41G2o+UX2JlfL/IAiGGNYGFSehkYe9VYZ5BcW55porDcn5zf9EAmGgglQxqlgNdRPpKl7D2SpWFTNxodIMgkkd/tAs3Ztuumm5JQgmDdTx6m1/CeI86ihP+66+ZlkmhhlgdPK4CrIcG5kkmIlhxhbtg+0MLM5HNAfDTwjpIOhQFE1DeqxxKlD4bmicSGaBEIuX9UHFyophAhgrHEudCptVToXtHCzkKmv/Z5+4TncdCbobIfGuvfbalGcNRS+11FLlL0HQOairs1hWx3K/YDVmMWYIyaM1/mf0UP+qx+3LVYnlmTGFYCauWYvt4xz+J7yDziWEdBBMwqi4cwxQlm2CWwVMSPs/W7T9tvDCCydhwk2EqFbxs3yLCcwqYljcMLchdxbtPAQY7iPBcKETaDEVeXGbbbZJ+TQIhoNsUfYhitWp6l4jg4SwUUNGjDwBnSsRQwVff3WselUdm10w8qih44NJmxDSQTBCUbSzRVuFz+LB/YOQ5gKiIrdQBSsI3zmrxRHhLNwqf/sbarQKGNFt4ldeESws2kEQjCQIZfWluo7BgRHBNqLY5ERCWL2ozjMXhssF1wv1pX34OM8zzzxpm7qXpTnXjyM5rnwQQjoIupps0dZQaAw0AiZxaTA0KCZ/GaZkfbGss8bD/9mizZ2Ej7ZGxn6EtwaIW0lYtIMg6CTUdwwLBHOOrMQqTASr28QlVxea4M2irA5TF3KdM1qnjlQ/2s/x3DT4KXPhcJ6gOwkhHQRBn6gaskVbQ8O6wlJjuL0vi7bYwiZBmhQjBJOGhbWG+4hjs0Vbo5MXRAiLdhAE7STXV+onHfkcyYUYNoFb/cO1gjsGNwyT9xgT/MYFw362MwowEKgDWZSN0IVRIOiLENJBELRMvUVbQ+Q7ccxSzSqtkbIKpP+FLqu3aGvwHCPer981fhovAtwkHII8LNpBEGTUE+oGEMe57jGSRhirM0zMY0Xme2ySn/8JYe5o6hv76OCbQ0IcC7PomHC/CFolhHQQBIOGhs8QKN/s3hZtDaKFBEyIJKot/6yB0wAS34ZQ+RkS5Ro/ViSNJ4uSRpFoJ7SDIBg5kCSsyT7gfqH+yBblbEU2uqUuES9ZJ1w9wXdZXUFUqztMTlX/ENTcMAjm6JgH7SaEdBAEwwYxbBa84VONIjR4hDTLtAaT+wjLEZ9F1myWJEtT5wk+lqDubdHWCGtQWasidFQQdA4kR3YZU5aVT98JYWWf0BUaTnQLHW5x86EuIJDta16GMp7Dx6lHHEcwB8FQE0I6CIKOJVu0Dd1qLDW8FixgneYmovFl0daoanw1qhpgK+sR3qxYLFr+GsLN0UvCoh0Eg4eyReQaQWJNVoa5TugsK8PmSNhuLgUrMnHMBYNYViaVa5Zmcy/sr0wTyTrGym8QdBIhpIMgmGTpy6KtwSakWbPMuiew/TUpkiuJKk+YKsPErNizzz57EuyGis3GB+tWWLSDYMIoezq4xLIyJWqPbVy4xK4niJVB2+2n/CmLylmeI2G7zi93LccSzspeTEIOJiVCSAdBMGIhsDXWrGMEMUsX8SyUlXja3EOyRTsvVOP/7G/JEkYUsKAR2Y4l1PleOl9YtIORCmmgg6mjam6DzigrsoVHzGPwv4gYOWScOQ7KBfGszNiHq5XyRxgrT8Qzi3JM7AtGEiGkgyDoWuot2lxG+GgS3VaGJAQIg0ceeSS5kli17NVXX00+2MQDlxHHsm7z3XaOeos2dxJiOyzaQSdCJMvr/rIqy8/kgDJACHPHYC3mQuU3/5vox8JsUrBjbbd0O3GsLHCZMpIT7hdBNxFCOgiCYAIQ2oaiWdIIYu4gLNascyY+schZqIbwICr6smizdLPMERjOQ6hYxAEhOILBRPMuz7Eec58gflmUdfJYilmRdRJz3pY3fX/xxRdTZ1AnkcsUC7I5B0S3jmQekQmCIIR0EARBy6g+CRLWONa6eou2yVEWdHj88cfTQjV+M7mKKPHd5CriJlu0ifY8/E3EONbvhs2DoC/kGfkF3I4IZp0zYlk+5GZBIOsMsiLr7Pnuf8fKjyzNOnms0vKcD8Hs2CAI+ieEdBAEwSBBrBA33D58WLD9JVKE+CPAF1xwwWS1FlFkgQUWSP6oBI7JWcQNkZ1XWSOWCHTCB2HRHvnIQ9ws5BuiWf7gc6yD9dprr6UOGh9+y1rz2Tdhj++/pp0VWZ7TMTOpVqfPdi5IzhH5JwgGTgjpIAiCYYJIYjkktolkAptlmygidggoftksiH4z5M6azX9bBATWbWHCDL8TRXlyF3Hlt7BoTxpkscxyzG2I5Vg+0GliXSaGjVboeFly33v2fp977rkUMs53eYCPMnci58u+ykR0EASDRwjpIAiCDiVbtP1VVRPPRDLLI1FNKJsE6X/ksH6slyKTsGgTZIQ4C2S2aPNzJbCItmDw8f7yqITJet6l9CeKCWI+8zpP3qd3ZYSCqPZuTYKVByyl73g++IRzjhjj+CAIho8Q0kEQBJMoqm/CilhmrTQJzNA/scaCzcppQhkRZnIYwc2CTbiJqW0Zdt9ZPVkwfXcMgc2VhACMEH+NodPCPUc6ex86LdLZe7E6nxEG6eodsBzrzBDP/tfpER2DWwbLM+HsfXifBHe4YARB5xJCOgiCYISSLdosnayZ9RZtYf2IZRZQkyMJNxPPWEm5h/Cp5avtOGI7I+JDN1q0c5g4wlj6eHaRW7jmcLVhRdYJ4dvuf2La/yzLoroIE0dY83nnjiENvZeIgBEEkzYhpIMgCLqUeou2iWzcBFizCWi+2AQg31uimojkZsBqSvyZ6MZ66nsOqUZQEo45+sOkZNF2rwQypIVnkh6EsnCGLPyELwu//1mRX3rppeQyI61YlKXBHHPMkSzTOhrSho96uF8EwcglhHQQBEHQJ9miDUKaBZYwJB6feOKJFHOYO0i2aLO0mhxpHzG1iXD/iyrhXKy6xCVByl2BVXYoyR0HQpfAd39cMDyHzoOOAus7qzPxzFrPykwkezaCWEQM2/maO4/nYeX3nMRzEATdRQjpIAiCoCWyMGXRJrS5O3AN4b5AkBKjhHiOJkKIzzTTTOkYwlV4NlEmRKmot2jbxqLdLO6HNZlg//Of/5yErW15Uh/xzC/Z/3yWWZQJfFZk7hisz1wwsuh3f/Bc4accBEFfhJAOgiAIBgWClEXXX+KZNZefMHFNxLIEE88Wp8kWbUKXpdpvvjcjqAny+++/P7lduBbXE9Zvbijf/OY30zW4q4iGYZIfse36XDXcY4jlIAiaJYR0EARBMGyYzMilIlu0he/jp237/PPPnwRvo7ByX3HFFcUiiyySLOBcMLhcEMlcMcL9IgiCdhNCOgiCIOgoWIqfeuqpYq655ko+yI1CkD/44IPFD3/4w3JLEATB4BJd8yAIgqCj4Kss9rJJf81g/7w4TRAEwVAQQjoIgiDoKEwKNBmw2age9q+PeR0EQTDYhJAOgiAIOgq+zCYANhuDWli+ZlxBgiAIBkoI6SAIgqCjMFFQPGqh8JrB/k8//XT5LQiCYPAJIR0EQRB0FJbMFleaZboZ7C+8XhAEwVARQjoIgiDoKPg6i/VsxcBmECd6zjnnLL8FQRAMPiGkgyAIgo5C1A4Ls+TlyRvF/s8//3z5LQiCYPAJIR0EQRB0FBZQIab9bQb7W0kxCIJgqAghHQRBEHQUXDumn376pl07PvvZzxazzjpr+S0IgmDwCSEdBEEQdBT/+te/0nLfonc0Ayv2L3/5y/JbEATB4BNCOgiCIOgo/u///q/48MMPi//3//5fuaUx7G+Z8CAIgqEihHQQBEHQUXDpmHfeeZsOZfelL32pWGyxxcpvQRAEg88nKlXK/4MgCIJg2Pn3v/+d3Dr4SjcTS5ol++9//3sS1EEQBENBCOkgCIIgCIIgaIFw7QiCIAiCIAiCFgghHQRBEARBEAQtEEI6CIIgCIIgCFogfKSDIAjahJX1/ud//qf43e9+V24JgqCT+MxnPlN885vfbGoSaxBMjBDSQdAgIgK88cYbqQKeYYYZyq3di6pDrN+XXnqpWHzxxcut3c0HH3xQnHvuuUlIizjRKBYgEW1isskmK7f0j/QX2YJ4//znP19u7R8RMYh9Ieb+8z//s9zaP/L/X/7yl+KrX/1quaV/6pf6bvYe//a3v6WVCpu5R3Gk//rXvw7JPeYIIUN5j955M6s9ukfpSDz+93//d7m1f+RHx33lK18pt/TPQO5RPv6v//qvQb9H11J/L7XUUsWKK65Ybu1ufv/73xdvv/12sfDCC5dbgmYJIR0EDaKyv+6661KjtMYaa5RbuxdiR8dizJgxxdFHH11u7W5+/vOfF8svv3z6zDHHHOXWiSMdrcZ31113Fdtuu225tX/kx2eeeSaJspVWWqnc2j/vv/9+ccsttxRLLrlkMc0005Rb+0fn4LLLLiv23HPPckv/fPTRR+keCc4VVlih3No/FlW5/fbb0z2yHjbKb37zm+Kqq64qdt9993JL/7g39yg9vbdGee+999I7W2KJJZq6x1/96lfF9ddfX+yyyy7llv4hGJ999tnif//3f4tll1223No/7777bnHnnXcWCyywQDHLLLOUW/uHsLr11luLHXfcsdzSPzpn7pFYXXrppcut/fOHP/yhePTRR4uZZpqpmHnmmcut/fPmm2+mZ9t+++3LLf3zpz/9qbjvvvuK7373u8X5559fbu1unnzyyeK2224rDj744HJL0DSEdBAE/VNtxCoPPfRQ5Yknnii3dDdVAVh55513Kpdeemm5JXj99dcrVQFdqQrVckv//Otf/6rce++9leWWW67c0hgffPBBZfTo0ZWDDjqo3NIYb731VmW99dZrOh9XRVJl7rnnLr81RlW0V04//fTKIYccUm5pDOm4wQYbVJ566qlyS2NURUFl/vnnL781RlW0V0477bTK4YcfXm5pjFdeeaWy8cYbV55++ulyS2M88sgjlYUWWqj81hhV0V4ZNWpU5aijjiq3NMYLL7xQWXfddSs333xzuaUx7r///sriiy9efmuMqmivnHLKKZVjjjmm3NIYr776amW33XarVIV7uaUx7r777kpVsJffGqPaQajsvPPOla233rrcElQ7JJWrr766/Ba0Qkw2DIIG+cQnPpGGHg1BBjUMkzYzjDvSkUd8PvnJT5ZbgiDoFHLZ/I//COmT4ZbEPSlonchNQdAghuDfeeedNFwa1Hx0Dee+/PLL5ZZAmvDd5CYQBEFnkX3vucgENcxzee2118pvQSuEkA6CBmHN+OIXv1h84QtfKLd0N9lCP+WUU5ZbArB4NTP5LAiCoUGdZUQxInb0YM7PFFNMUX4LWiGEdBA0iOFAs/rDlaEHgrGZWfMjnTx0HK4dQdB5qMPVWVE+e2AMaSZaUPBxQkh3GEIIvfrqq2l2fLcjlNKll15avPDCC+WW4cWwoFBBZpkHNTcGEQ9E7ghqSBPhzWLoOAg6D3W4SDLcr4IaQlq+9dZb5begFUJIt4gGUxip008//WOfM888s3jwwQfLPRuHiH7llVeKY445pjjuuOPKrY2h4a6/h3POOSdVGs8//3y5x/AjLNLjjz8+3n3mz1lnnVU8/PDD5Z61GKHCWO2///7FAw88UG4dXlgbDYM1Ex94JCM9DJGGq8v4sHqFxSsIOo88YhSTDXtgoY86fGBEbhoAxB4nfQswXHDBBcky9/rrrxc33HBD8eMf/7hpMU2ciwnL6tkoxPevf/3rYvTo0cWFF16Y7sGHICdQzz777HLP4Sd3PliY99prr5Q+7lUaigd6+OGHp3iW0AkwqY91r1NQAX/rW98qpp566nJLd6NR4jPeaLzkbkCa8MHU4QqCoLPIHf9mFn4Z6XDNaybGePBxQki3iAbzG9/4RnHyyScXiy66aFo44LTTTksfgc2fe+654qc//Wm5d2MQagLnb7TRRuWW/iHmTzjhhOLyyy9P1833wKptcQhuIp2Cnu/KK6+c7o3QsLBDfZpZ8OGII45I+/p9iy22aGr1r8GGuLfgQyz/XCN3/KxsGNSQJhG1Iwg6k7zSY7he9WA11k7SCZMiIaQHASJbj3fyyScvt9QaWCKM5diH60Um+0Xn7Qp6I2RXECs07bTTTsWaa65Z/lIToqecckqx8cYbp++ub7UwLhT33HNPcj9h/c3b832xrgtpBpXOE088kbY7LluLWYmtDmV1NKt05eOs9NUKOhDTTjtt8aUvfanP2dTukV9y/XUIFd/PO++8cddVOVp50Hbp+OKLL6bt7cJ98NuOSrgHnQt+0kEPyqV0CYKgs1CHK5vKaFBDO89vPGidENJtQKHki0zAnXHGGUlgrrfeesUGG2yQfld4iegrr7wyuX6Iu3viiSem/bKI/slPfpJ+87/lUhuBoCVuWXpXW221cmsPxPxWW22V/if+TjrppLR0Lt9j1xIT2ZKplnj2nWXRffzsZz9Lhevpp59Oottvnu+QQw5JS+k+9thjxUEHHZQ+zuU4wvXaa69N12qE7AMtzXy4xrA+97W0r/RT0PlK77vvvmk5ZfdnOdr83fPdfPPNablTnQvLC7PUtyru+4LgtxSwkYighigmMSzYQ7h2BEHnwlCjzgrXjh6+/OUvFzPOOGP5LWiFENJtgNAzPEJQ7rHHHsm3lzV47rnnTr8TfUTzRRddVMw000wp0yrQhx56aBLDV1xxRbLq8Wkm/hq1ZhHhb7/9dmq860OQuR4BnEUqkcsdgeA0yYJP66hRo4rNNtssTfDzf74vFQx3FVZqnQJi2m/TTTddsvCKouFZ//znPydxK2yO/ZdYYol0zUbxjO4ndx4I9a9//et9+kS752mmmabYe++9yy1F8nPjIgLpL835WBPo7ldcTL7qLOrtwnW4MjQ6YtANSG+dsaCGPCJvK4NBEHQW2kx1VowY9cAIpU0PWieEdBtgqVxqqaWSePaXpbQ+nIxCaxtBSDgSv8sss0wSn4TjTTfdVKy11lppXwJ7xRVXTP/3BwFNUKoc6icoZmH50EMPJT/kp556Km1jvXX+eeaZJ+3nvohjFjT39Ytf/KKYd955k4sI1wmWZwLfbyzq22yzTbI+LrvsssUiiyxSzDnnnMmP2X00G4eSxc6Ewxy147DDDkv3fMABB6T0aQbPz/XDfeoAvPnmm8lKzxrPXaRdSEPpEa4MPci/UQmPj/wYQjoIOg9lU50VQroHQtrqhkHrhJBuI6y5onUorCzLrJcZInq++eYbJxxPPfXUYo011kj7EoB9+Qb3BwFP+Oph109sJCK5ley3334pVBtxyge5L9wXa3P9fZns6BwE9vrrrz/uN64hM888c3lk+3APImEQ6lwxHnnkkfKX5rBQis6CezWB0XO3M9C8+/za174Wq0DV8dnPfjbln6CGTqWyHEPHQdB5aDMZcbRvQQ3GuO985zvlt6AVQki3EUJrwQUXTO4dV199dXKrIKazWOVfnOM66xUTv36bYYYZ0v72zcJamDiROCaGBlu0kMUWWyxNHuQi0gwqFeHchKDLMZz1TrlvuI/pp58++RqzdvvOKn3XXXel/dqN67LMEyJ8tnqTre/ZKszix5pu8p/jHM+9JaeZ9OXWIbReu3Bt1/MJarDshKvL+MgnyksQBJ2FsqnOivLZg7Yy6vCBEUK6RRRIYlc0C77RBLKJevyGTTRcffXVk7sCC6+JdKusskqyZgrvRmCLNvG9730vWa4Ib3GU7SvuM/FHGHK1cA2+yn2JZOJyqqmmSr7Bwsr5m/2iHWMy36yzzpoEKD9W52C95jtMHBPi3Eu4ephI6Dj3ajKd82655ZbJf9nESEKdYOXSYdKfCZNcMGzLExDzdwJWWvRekZD49ZsoI+6jfrKhDx9y1vCFF144idWxY8em5zf5UhpPOeWUyb+bWJZO999/f6oU+X+LkMKVw7mdK0/eFE6wXbiWmN2//e1vyy3djTKg89cpK092AtJE2Y1Z8EHQeWiDRKVSRoMaXPNM0A9aJ4T0AFAY+ULPNddcxWyzzZbiNuvdGTYyMY6rQvbZNQGO2weRSuCZaLf11lunfblP7Lrrrmlf4nmdddZJ4pprBkEpkwvrVu8qkmFVXmihhZIId5xz+7gXvcx99tknWWoJV5Zc1/S/8xLiolAceeSRSXA7Tji7TTfdNN0XX20+1p6T1dow/uKLL54KHvEtfrbIH5YYNTSUvxPthLYoGvUQGX6zD5HuHvL9Eqe77LJLuhf3y2JA7PMdNwnR5MbsuqHzIZ10RKSbdOW7veOOO6bz5udwj+0cssoW/FiQpUYeJeArH/QQUTuCoDNhPFJnhetVD9pb+iUYAFVxE3QwVRFbOf300yunnHJKpSpCy62dS7XHX6mK6Mro0aMrY8aMKbeODKodkMqTTz5Zef7558st3c2///3vSrWzU7nhhhvKLUG1A1updiwqt99+e7mlf+Sre++9t7LccsuVWxqj2qFN5eyggw4qtzRGtfNfWW+99SpPPPFEuaUxnn322crcc89dfmuM999/P9VfhxxySLmlMaqd4coGG2xQeeqpp8otjaF8zj///OW3xvjjH/9YOe200yqHH354uaUxXnnllcrGG29cefrpp8stjfHII49UFlpoofJbY7z33nuVUaNGVY466qhyS2O88MILlXXXXbdy8803l1sa4/77768svvji5bfGePfdd1M7dcwxx5RbGuPVV1+t7LbbbpVbb7213NIYd999d2XppZcuvzXGL37xi3StbbfdttwS/OpXv2o67YPxCYt0h8Myy6LN6t1Jq/xNiGqeStZjFmHuLCMJrh2s6bGyYQ3v2jApt5ughjQx4hMrGwZB56EON1Ibrh09iNjRzrlE3UgI6Q5H1A1uG8LqTQoYOuPjfPzxx48X23okYGIoX+yR9lytwrWDC8O3v/3tcksAZYB7RxAEnYU6XJsaUTt6sEANF8+gdUJIB0GDEI7iUvOxC2rpwdcwwgH2IE0I6Wiog6DzIKR1cs13CWroWDAQBa0TQjoIGsSwoEmiwgAGNTcGE02fe+65cksgTQwbR9SOIOg8ImrHxxEZSyjZoHVCSAdBg7A26r37BDVYXw0NBj3IJyxfQRB0Fsoma3SUzx6MnkUdPjAiNwVBg0T4u/HRKH3xi1+M8Hd1SBPuLkJFBkHQWUT4u48T4e8GTgjpoCsxBC+ygmG+Rj+ikYinLXZ4X79320dc83fffTctyNPX7934yREBImpHEHQe2bVDOe1ddrv1IxIV97y+fuvWT7OrF3+iKigq5f9B0DUQO1ZhbGZFJ4vtCPVmKGz22Wcvt3YvQjNaYOepp55KK2sGtVXC7rnnnqYi7WjcLWBkaf7jjjuu3No/xMDdd9+drrn55puXW/tH58cKoBZwslBUo+hAisZj1dBGsQiU/OFemwmH+Yc//KG45ZZbiqWXXjqNAjWKlUetfGohqkZxb+5R52ellVYqt/aPBaNuv/32dI/TTDNNubV/LCZ1zTXXpMWuGkXj/vTTT6d6a4UVVii39o9QnbfddltavKoZq6PVSi+88MLilFNOKbf0jzBq9957b7rHDTbYoNzaP96ZutgqtM2sRPvss88Wl1xySVp5t1HMb/FMDz30ULHaaquVW7sbaSL83XLLLVdu6W6070ZZm2nTQkgHXYlG87LLLkvW1EYhHIkW/nURAq9m1ddzJ3oiBF4NeURIQKt0Npom0pFQsrqnFTobhQA3UUjc6maEnHem8ZxqqqnSaqGNYgIlMW2Z/omhbGmYpcPMM8+cOqBi4etg8MUk6myHyap33XVXErP121F/HL72ta8Va6yxRhoVItggtj5B1MhzOJ/49joSiy22WLl1cHFNq8wSwd///veLGWecsfylByva6jRIAxFw3Nt7771XzD333OUe/eOdmjAmbaw+O9BwZkabWCqteNsonlV+VAbkrUaRX9QhIiJ9+ctfLrf2j3tstsw45s4770zCvZm8P5KR73SCmqlDRjKiuqiL1ltvvXJL/4SQDoIGYWl58MEHk3/dUDXEnYwGU2N76623Fttuu225tbvh/mNpfGKmWxsmFteDDz44Wbg222yzZLkdNWpUEuGEEgFz5JFHJn9ylsErr7wyNV7mHmyzzTbjQnEpb0888USygrPY+2333XdP24455phkRd51112LHXfcsSEB5nzO4z5Y49sB8UgEakb7Eq8E7v3331+cfvrpxfrrr19svPHG5S81pM0FF1yQrKs6CiYyE5TEjeduFPsThxdddFGx1157Fcsss0z5S1APIc3aru5SRoMidXoff/zxVFaD1ggf6SBoEI0lCxrrYdAT6o2QCGrUW4m7EYJOoywNMiyuOqAnn3xystQ///zzySpsu04HgXnggQemtHvkkUfKo4rUYV1wwQWLnXbaKQ217rfffuO26bix+DuuUSumY+edd962iWh4zuuvv7549dVXyy3jQxiz4Pcl2ri93HfffckizxXljDPOKHbbbbdkHWw2fCJLP7eIZqzY3QgBrf4mqIMaRgSUxaB1PvnjKuX/QRBMhCwcJ5tssmLKKacst3Y3Ymv7NONrO5LRUMsjRF4eOpZvbB/pIbdYZ1l7H3300WL66adP4o6w40fPdcEojjQxL4H/OPeFa6+9Ngll26Ubn+8VV1yxPGNP7HbWZ4I7b+Py8cADDyQrNQgB1liuWv5n3X7ssceSW4iOnnsiXIlWKMME/XXXXVc8+eST6cNXd4YZZihef/31ZCVnvfbuuKgQ/CyZ3qHf7GvEgRX4vPPOS/sR9CzQXMZYmD33d7/73STcHCtaRH2EG+fgh6xjkIeRWaPnn3/+tC+LPX9v7hrul7i+4oorkvBxT1dffXXx8MMPp1Eh7g0EuOefbrrpUv57++230/Gex/7OSfDfcccdqaMnnb7+9a+n645kvBtpCeVQ/hFtqBuevRGUW/laXg1aIyzSQdAgKmQNpQY/qKFRIlCCGhpqgod1VX5h+eKKQAiOdDwrP91FFlmk3FKDy8Lyyy9fHHbYYUnELbvssknEcIMRjowAFVrSJB9uIb2Rx2w/88wz08dkR+5EGVZh4pYl3Ieg5kNNNJqIZhInMUmQE+7uwTsinu1PjHK9ILZdhxAmormdnHPOOUkEE+V77713+s12kzVZ1XUGPAcxqxNh8qHJffZxH/WW+d4Q2DoEvTuhXFtMYCSMb7jhhjQBlaXf/Az+vXyuPZ9OAUv/ueeem65fj/u66qqr0nNwLSH27eN4x9x4443p3CMdnRmdKe9G2cwd3ajDeyCkow4fGCGkg6BBNOisSCa4BLWOBfHEshfU0ECzuIqWQLAQfieccEIS04TTSPxohD23ssF9ovfkL0KZeCYqCdNmJqJBPnMdotBH+roWlEkWW8KaHzbRKTrFmDFjiiWXXDJZmOeaa67kk83SnSM1uE+Cn6/1JptsUqy99trFVlttlfIy8cXNgisJwa0T5HedI5MbDznkkNQ5IGxXX331ZFHmX+oZv/GNb6RoHNNOO20qG70Fbm90JFhHe6NT4b7333//9Ays+6690UYbpUmLXEIOOOCA5C7Dmk1oZ9wnv1dCWlo4P4GvY8EKbbTgO9/5zrgoHtKw9zsdKR8COpdB6SENTLTt7710E/KxchW0Tkw2DIIGMRxKEJkYpfHsdlh3WOVYvDbccMNya3fDh57PrElkxB1LJj9ZAoggGomINMGCylJMALIue25iky8z4czFgFsDFw9pRATqbBCy3BXAkkvwEdsZAp1oPOuss5IbRt5mX+KY5Zd11rVZm4nILDJ/9rOfFYcffnix6aabJos4wcAdwt999903jS6Jn8tFZIkllkhD28LSsQTzWWZpJr6EvBTOzbNw8SDQjjrqqHRe7h35/4UXXji5VqgjROlgFSZ0pY97kQ71kw2JF/dJjG+55Zbl1pplX+dABBNpxaLONWPRRRdN98ZF4+ijj06dhfrIE0Qjy7P9pJFn9Nzgiub/7CYjL/Ldds/eA4v+SEQ5lG9Y/r0rnZ2FFlooRSMRmSGo5RvlYK211iq3BM0SFukgaBB+dhq0WCK8h7xSWFCDryFrJ7HlrzCJxJ0OB0vnSPxkFw2izmgNaygRScT4EG/EDOGy3XbbJSsv9wTuHT6EKvHI0kzQNgPR7rrOyX2DXYiY5yc8MbK7CGE8zzzzJFHpu7Lt/j2XjqLzNxrGkLVXXGN/Wa1ZfScGcctvnJuF9EAOY8fdRL6Rf8Ss545C8LhX+crKmTkGvhGBfDzcM19rYpFFW9zkLbbYIlmmWaNZz70nQhyG9nu/05Hy0fHgUy5PeP7s2hF1eA/SJpYIHxhhkQ6CBtHIsYSphOsnRHUrWYywZmmwg5q/Luur8GMacP6ZhBE3gx/96EflXiMbIpp/MKHIEs/axYJqEp3OKGsrf2MTAlntjWgQvkTP9ttvPy6MHIFH1LJQsxofdNBBKY60bVwvHCtEHBcIPs7cG+abb75UTsVrlj+5elhYQTQMVkmi0j2YpEhEE6hbb711EqPE/Kqrrpqs5NweWNSdgwVTNBHXECXEiBR3AQvMrLnmmmnxHVZnUTOcj48zsctazlLPEs+PmSAXmq4+TJ7yI22IZsdrjglhz5EXJ/G8rO8Wi5GeBKI8xuptH/fDpYRAZJnnsmLRFtZpgpt49szSWH50Hzo/znPaaaela4xUuHIce+yxyQAiHKN3YRImQd3M4jsjGe5MRnWUkaA1ImpHEDSIyldjr/dOBAS1zoU0qY9G0M0QRAQKNwHD5zkkGWHVzAp9kzLEIAHKlcEz85EmSk3u4x7F6qxjIU34/epo6HRwcahfAERasmab7Oc8zsk/2DZWbGKZ2BZazoQ95+EKYQjfuQh2v7s+sc1SbBsruG0EPwFsOxHunRn6d6+u6V5dj4uFzoDnIXLdt5EH5/B+fWd59zsrNMs4UctP2jMQ1vKEZ3XPOU42RONgceZu4T4cp8NRH6feOWx3bh/i2DnyMSyKOm4Wm/EcrNFcz1w/pwnxTtT7nYg2YqKD0Z/lfiTgfXPNka7elU4TY0hfcb+7EXnCiE4zi+8E4xMW6SBokGwhM4zdzGpaIxVVBwusUF+xvGwNjTQ/WY0S4RQEA4Xg5+pBLBPJQevosOlwMIqEcKzBzUcHU+c2aI3wkQ6CBmERYw2LGd81CGnWLta6oAbLId9VFr8gGAhGekx+NHmVa0KI6IFjlEH9LXJHUIMxxAhP0DohpIOgCXJg/6CG9BjpC400S+SRoB1wm+LXbUGZcJ1qH8pnlNEeIj0GTvhIB0GDsMCyOGafz25HevDf9Bmpod2axaiFPML/ki9rELSKaDgmDvIB7yvWdNA8XDqUUfNcog6vwUqPbvCXHyzClBQEDaISNmlIHNqgBqtZDJP2oFMhLq90CYKgsyCi1d9Rh/dgXkcsMjYwQkgHQYOwwBJIIZJ6IBzDH7gHnS2z4KVLEASdhfJpxCjq8B5MoldnBa0TQjoIGkToK0P2wlwFNQyRxuz3HsT0FeIsFjgIgs5DqEAxt6MO74GrovCRQeuEkA6CBgnXjo8Trh3jE64dQdC5hGvHxwnXjoETQjoIGiSHewtXhhp58qU4t0ENQjovrBEEQWeRXdGsYhnUEFtbnRW0TgjpIGgQrh1WFosVsWoImSSagJX7ghpWTLO8dERZCILOw8qG6m+rXwY1LBxldc2gdUJIB0GDZAtsDhcU1IZKDQ0GNbj/sPBIlyAIOgvlU/0ddXgPrPTqrKB1QkgHQYOohN99991wZSjRsSCiLS8b1NBAv/3229G5CIIORIQKC9xEHd4Dd8W33nqr/Ba0QgjpIGiQ7NrxrW99q9zS3WTXjnnmmafcEoRrRxB0Ltm1I+rwHrh2zDHHHOW3oBVCSAdBk7DEBsHEiDwSBMGkQiwRPjBCSAdBg/B7FepNeLOgJhbNgH/xxRfLLQEf+tdffz0WOAiCDoTrlfo7wr318OGHHxavvPJK+S1oha4U0gTRLbfcUjz88MPlluYhIt55553i/PPP76hwaHzAPNujjz5abhlcTFR4+umni6uvvrrc0h48xwMPPFDcdddd5ZbhJ7syfOELXyi3dDfSwwIkX/va18otAfcfQ6XSJQiCzkL5tFhSLJjUA3e0ySefvPwWtMInqoJw2Mcg//znPxeXX355+l/jbKWd9dZbL303wctv4j4qBKuttlrx9a9/Pf3WKsTf2WefnQTAuuuuW25tHEkmoPvhhx9enHfeecXLL7+cfGd74zq33XZbEtyf+tSniiWXXLL46KOPimmnnXZQxJjr3XPPPcXee+9dLLvsssVJJ51U/jJ4ELx33HFH8cILLxT7779/uXXgsOxdddVVaTbxVlttVW5tH+778ccfL371q1+VW/pHB8xElUUWWaRYaKGFyq3di7LJQn/xxRenPB3U8u0vfvGL5IcZjXUQdBYs0jlm8tRTT53+djsMgZ/5zGeKTTbZpPiP/xg5tlXtk9GHp556qqnJ37TadNNNVyywwALllv7pCCFtBu0hhxxS3HrrrWlIdNdddy0OPfTQ9Btx6DfCd8MNNyx23333Yvrpp0+/NQoBdOeddxYrrrhiuWVgSDIvaLvttkvCtS8h7SV6gT/+8Y+Lb3/72ymDEhust8ccc0yfwnugqCR+9rOfFUcddVSxxhprDImQbhfu/f777y+WW265csvgQqBfdNFFxRNPPFFu6R8i6aWXXiq22GKLlEe7ndwZ2XbbbYvvfe975dbuRr4SxUSZ/9KXvlRuDYKgE1CH0xva58FogydFrNbLeHnmmWeOqM4/8XzzzTendn7KKacst/aP0UTGMh2LRukIIQ1i98ADD0xCkAW3Hg02C/U111xTbmkcj/faa68V22+/fXHfffeVWweO+yWiCda+hLQCu88++6SOwBlnnJGe4dJLLy1++tOfFhdeeOGgFWIdEVb2WWaZZZIR0iq1n//858XWW29dPPjgg+XWwcU1VajNuOUYFTn66KOTtfG0004rt3YvOj933313sddeexXXXnttubW7kZ/k4fnmm6+pyjsIgsGHuNLWqP+V0aBIuuiKK65I+mQk1VlGHsaOHZv0384771xu7R9GTy6czbgsdoyQzoJ3scUWSwJ1zjnnHLf9zTffTBOafvjDH47bxupz7733jnMFIR4VDn7PBI+PRu0b3/hGauRvv/324rDDDiuWXnrpZC3iNkBsuo7zcS+R6MguJBKSI/6VV16Ztktgoa0WXnjhfoX0P//5z2LTTTdNwwRHHnlkGiogqmXaueaaKwltvSX3/5WvfKVYa621kruI+9Ij2njjjdN9zzTTTOk41m3bN99883R+13/uuefSdufgl+kcWUjPOOOMqUeVj1t77bWLz33uc2mShbSYYYYZUhpa0WjBBRdM2/lWw/6rrLJKen7Xef7559Nw9RJLLJF8of/zP/+zWGqppZKF3b3xx/a8rMn+6gHWIw2kmzBpjvde3PMUU0xRrL766sWrr76aRhzGjBlTnHrqqel+3D+RJm1YO70jPefcmXKP7kG6e+9cDKSt++ZqwjLo2dppKRVv86CDDkqWRu+029E5JBq59LBMBzWLtPrgu9/9bqqXgiDoHLRPRpO1J82ObI9UbrrppuKUU04ZkUKanrL2AzfcweSTP+Z70AEQVpNNNlnxyCOPpIaIwAKRdMMNNxTLL7988dnPfnaciPby7cd6TYBZpljC7bfffuk3Yo84dF6Cm/WRQz1hSlzusssuSWR///vfT2KZ1dh2Yo2AJTrnnXfeJHZ/8pOfJEH50EMPpQlwxLPzE5f8t3fcccc+G03+0GeddVY6P99ay5IS7vyR3NsFF1yQhKOYlnya3f8ee+yRzs3a5x758Gqc+SCfc845KR08xzPPPJN8Uz3/r3/96/SbNHPf7ikHnNcBUUD0vv127LHHJhEorYlPfwnmk08+OaWn++QG415mnnnmdH1uNsSx44l3v+t4LL744sk1grgUqWCdddZJPf599903vTf3xfou/XPn4+CDD07v0LWMPqy88srpXvWI3Q+/Ne9FgPgDDjggpQOBLi2llfzh2jpMOljuUaeEu4yPOKE6ZO7LPquuumoS3e1AJXzdddelDtVKK61Ubu1evE/vQH7g3hHULF6PPfZYysMRSzoIOgttqbaFUYRBLSiShV6dxRA3klw7aAbRSBgXGd0Gk47yLCdQNMgso1YHA+sly1eeVarxvuSSS5LAZeEkoAlVbgwEGSGssBBsRCyT/g9+8INiqqmmSmLZMQoSgQaCjzWNQDJc7xhCEASf6x1xxBFpO5HLAuca/cEKu9FGG6XnkVF32GGH1OvTQ/Kc2fWCpdYzEPx6g8sss0wStZ6fcPNMLLTujeBmBXfv7ocVmiV39OjRSTASmHDf/s/HeWadAOlC+LC48wFynE4By6/f8/PzQz/33HNTxAxWcj149yJjSkMjA/zZXcf9vf/+++m60NmRXs7Nl5hI32mnnYo111wzncPEQdfgx+18fI5N3JNWJmC6B5ZvHYTsdpEt8qzR0owvlwmV7iFPSPRO7ec4714nhJCuv7eB4nldwyeoofz4BDWkhYo78kgQdB7Kp/ZCWxQE7aLjhDTrI4F42WWXpUxvuH7++ecv9+gRvgrDs88+myyuxCAxylrLSkqkTiicC4HLgpx/dz6Ci0uJbX43qZFPtf832GCDFG2D0Gx2+JollKgkGjfbbLNkJd1zzz2TKwThzGrFVYPA1kP+5S9/mVxAHOf6fidAuaPYP9+zjgVB7XnBwp0FM9w3Meo4aco9grBm7dWx8Dv3EhDlOi6LLrpoSnfWcOeVhtKFawRLN79gFmL3ka3veV/W5oxtru1ZPJeOgqF/1ySYiWvWax2hCVmKWZW5pxg9AIuz6CezzjprcidxDZ0E55M/WPp1VPSm3aN0GgxroLR03ojGUENe8A69j6CG9OCWFHkkCDoPdRWjmk8QtIuOi3XCWsq3mKWRJZRg7D0pgKBZYYUVkjXWh4VyINEeiMls/ayHyOZCwTpLsPHlbRSWbL7InofQZIXlp0PMcukAcckXm8hlFTZEztWhEYjLZkK6TAy9c2mdkb5EbLbaN4vzsVzzU8++SdKSq4dwgUQ0V5VGz88SrONUf4/Sjo9bq/fYCu7D9XRkglp6eK8+QQ3l3ijOUObLIAgaQ11lxMgnCNpFxwlpIs6EMb65rKy9Y0azghFQLMTZ/YMQ5WM7IbJ1SCEi4OpxPZZc1u18PvvxxSWY3AMfbfckDB8ICP7RE0NDyr3BxDcQ1CzrBGq2xGarNKsz4ckvmUW6P4hIMQ6vv/76ckvN/aGVRVjcl+fnI8XNAsQAVwnW/WYh8I0m6ESwDpsM6P1IXwKakGZV5r7CAu5arNf8r+E58n1kWBHmmGOOtD2PCthPHhls36d6vHfPFyKpB+8vhHQP0oOrWXS2gqDzUD4ZoEJIB+2kYyYbZrLrgEgRJriZQFY/DON3rgomFPI9ZqW0r+HUHGHDhDlizcx5ZKEt2gLhyMXixhtvTALNZDUuA4S5iXTOxwrN/cBERBMZc+B2Fml+w6JNgEh2Lr7NJhFyScgosIQjSze/ZPGjnddEOBb3LJgJeccTlsK/uR+NsPv1jES3ffkIE85+I8Z1Jkw2hHO7d1ZbopTwZxUmYnUO+BazkhGuXCSefPLJdE3ilFuICYec8nUe+BTnc4mT7ZlFM9FxkA7u1+RFz+G9EP/Oz2+c+4f9+Ce7luu7b/GhiV73xKfaJA/bpZ33KT0dy1LPp5rvtDTzHISrCCPu1bPxi/a7e5S2W265ZbJ8Swvp4LncFz96z6Mj5tgJuZE0g3vxLHy5hyredScjj5sgajLpNttsU27tbqSJfMndKHcOgyDoDHT61ePm8gx0YbeRQkw2HDgdJ6RBrJlYx/Lae1U7woug85EBfv/73ydxzKeYcCIANWJEcl6ZRuYQAoXYIw4JP+fX0PlLBLPKsnY6H3EoAgVBRmTm67gvItYLsrgLH2LH6eHysVY4eyMaBwHseCKViDahMON5+N2axLjbbrulc7C2ihyS79F9EMREr+86Cc5L0BGjzq2zwP+Z0HeO7CdMZEoTwlZ6Sgf+0Z6BX7TzEbLEJmu9cxECfLt1aPigO4aYJYRZ0Ilr351XOttOCHsPhES+Z+fy8Ts/c2kl4kpOC1FRVGys/cS17XzFpb2CnZ/DR6fG+xTtw34Kh0VRHCcCinTwHt2TjpH09N21TayUdgPFuXREdJi4FnU73rXODbekENI15BGjOcpJ+EkHQWdBRDO0aWOzgazbCSE9cDomjnS3QkjKyKyvFnAJOhdWfaMGRkT4zXc7GiWjMhZS6u0y1a3ohJ9//vkpso1RsiAIOgd1OCMLI0Bel6LbiTjSA2fkLKw+iaFHLN4zn2GTDFmYg87GiAT3ICMBQW00hXXeqERQQ3oYtQprdBB0Hlz8jJaGNTpoJyGkhwk9Ym4TfH35anFzCDofojGEYw86Fz5BDWnBpSrySBB0HsonN792uPoFQSZawGGC5Up8aaH7+AQHnQ8vKD7c/M6DGhEOcHy4u5iI21c4zSAIhhf1lTk1PkHQLkJIB0GDZFeGdkQAGSmERXp8TLg1sTfySBB0Hsont6twvQraSbSAQdAEBFKIpB40TD5BDWlhMmrkkSDoPHT6Q0gH7SaEdDBkiFBidUPxwQczID5XAzOzhWVrJ1w7hDoUVieoIa3DtaMHaSGWeuSRIOg8TPIXzcEnCNpFCOmgbWShfM4556TwcGJhExZ5NcLsY2yCJV/SwUBF6XpWoRQRpd2wOIYrQw/cXXyCGtLCRKbII0HQeSifRotiMnDQTqK2D9qGxShGjRpV3HLLLWnlQlZhYvbqq69OvxOhFn4Rs5If6WBAzFuwxeI77YY4skiNEHhB+Iz3xac//elittlmS5E7giDoLNRVFg+z2FkQtIsQ0kFbIGAtA26Zb0L5rLPOSisPsj4PJSpKqw4uvPDC5Zb2kS3qEZGhhvSIqB3jY6Tl9ddfH1TXpSAIWkNdZYGOiNoRtJMQ0kFbyJZgrhXPP/98st5avvu0004rFlxwwbSP2NlCg1188cXpOwgPC9NwBckfPtT8TPmxjRkzpnjnnXeKm2++OYn0e+65Jx2Xz1V/jOWqBxPCUUUcwrEH790nqCEtdLSUgyAIOgvl8x//+Ef6BEG7CCEdtAXC+Tvf+U4x33zzFbvttlsSvSb7Gfpfe+21UwXGYn300UcXe+yxRzqGIL3//vuTEH7iiSeSS8iOO+6YXEF+97vfFaeeemqx/fbbF6effnraz+98n//whz+kivAnP/lJEtgPP/xw2peYHkw8Y6xs2EP4G34c6RErGwZBZ6KuipUNg3YTQjpoC0TmNNNMUxxxxBHFEkssUey5557FfvvtN85SzJprIZN6qzGf6ksuuSTtTxQfd9xxxbTTTlusu+66yZf6lVdeSZbn3/zmN8W2226bzm0bazURJ8wYN5IzzjijWGmllYpbb721PPPg4BkIePcd1NKD5dU7CmpID0PHkUeCoPNQV3344YfpEwTtIoR00DY+9alPFYsttljyj95uu+2KWWedtdh7773TBEQCdJZZZik22WSTcu+aRdOkrPfffz8J8SmmmCJZfFkNPve5zxUHHHBA8dnPfjb5Wk8//fTjTVD0+8EHH1x84xvfKK655ppkwR5sspAerIgjkyIhpMdHehgxiTwSBJ2H8mmey5///OdySxAMnBDSQVvgusES9/LLLyfxe8wxxyRBvdFGGxU//elPk1W5NyIcrLHGGsW9996b3Dt+9rOfJSGdfaonhklu3DouvPDC4tFHHx10/2gQ/qJ2RESGHiJqx/jI0zqQ4f4TBJ2H+srIaUTtCNpJCOmgLRDSRPTxxx+fLHJQaRHSBCiB0RsWXiywwALFk08+maId7L///sm9Y2I4zsTGAw88sHjmmWfS34033jjdw3vvvTeoUTVYX8MC24N3kd9jUCsHrNH+BkHQWairGGF8gqBdfKKasaIVDAaMITMRNfgsr7LKKklE2/bss8+miVcnnHBC8eqrryahbaGWM888s/jhD39YHH744Sm+dL14JrqFsOMSYhLhPvvsU2y++ebFVVddldw59tprr2K55ZYrtthii2LLLbdMVuyXXnopWai5krAa87lWWR511FHF0ksvXZ55YHzwwQfpes7rnrodk0V1gPi5S/+gSJFmzj///JS3Z5xxxnJrEASdgDrc+gaMIcpoUBQ33XRTceihh6a2dbLJJiu3Tvpw4XnooYeSqygdMJiEkA7agorprbfeSguhcLVgXQYRffLJJydRbXsOfWf7kUcemcSyyYMZ2dG+P/rRj5JAA1cRonn06NHjvm+99dbFbbfdlq7Dv1oFwO+NH7Zhddci0Oedd960bzsQG1g4v/vuuy9FZuh2vCuVFd94LjZBrfLWofze976XogMEQdA5qMMZdIwYKaNBkaJeMWgxZo2kCEx0hPe8+OKLp5HxwSSEdDAsyOBvv/12CocnVF7GsPjtt9+e/NjmmWeecmtnwAJrxUYi/bvf/W65tXtRdWiYVFibbbZZubW7kR6WqJ9zzjnT5NkgCDqHjz76KLU72h9lNCiKn//858kqPRLbNAEKvOfBnrMSQjoYFliwrXq4zTbbpFjRGRUcH2fh8zoNIc1YwbmerLjiiuXWoUVH47HHHiveeOONckvNur/++uuX34YO79BowpVXXpl824cTeYZrDyFr8uPss8+eRiOGGhFoLDAkHON0001Xbg0mRbgB6NT//e9/T9+Nei211FIp7GYwaWLUUkdXO6OMDhfqK+2fEVVLli+yyCJpNLe/+UGDgQXUTPi3/kPQGp/8cZXy/yAYMrhjaJC4aRCGlmz10XjxXRPWrtNQ+bo/wlXlNxzwz77jjjtSzG0TLt3PI488khbCGQ4LqM6Fexgu6w4xL2IL/3lDlMIg+m7Vy9lmmy35zw8lRi34SVucKCJ3TNoQNqIJnX322WnOhxj2OmnyVTBpYvRMZ5sxZLjqcPfw4osvprkU6isfq/cS+cORt6SHT+Tr1gkhHQwbfGu5b6y++urjPiuvvHJHimgQ0ioc4n/yyScvtw4tfNi4vdx5551pYqdoJSxmhOPCCy9c7jV0EPbSZLisr0T8SSedlCzjJsyIU866wwVHOMZGQim2E8KetenrX/96yifBpIv3Z2jYKIPJy0S0ESn1VDBponwa1dMxGi7XK+4l3AMZQnTSjHQwBPDZtl7CUMMYIk10/oPWiPB3QdAg2frZV0zsocI9CC+o8ptrrrmSkCWihyO2Na8wq1UaohwOVP6iwrz55ptJRH/7299O2y3W8/3vfz+FRhxq3BPL5WCGYAyGBu+QtZBwthCTcj/UIxxBe1Ffeo/DWYcbjWURV1cwAIjus8ceewybRVhHMaIuDYwQ0kEwCUFAP/DAA6kyPu+889IiNmJnCwc4HBDTwzXNwlDoDTfckHzss4iGzobfvva1r5VbhpaYdjIykIfuv//+NBlLOSO+1llnnfLXYFJmOMuokQ5zOBg/RDvi0mhkdrii/AxnHT5SCCEdBA0inB63iuEMa8Yydvfdd6dhOJNmWDTE/xyuYTl+wBqFoYabDR9WlpTeYaxYEk2eEfZoqDH8LzQiP/pg0kVnzNC7OOlGPQzBr7322mmkI5h04Rqn/p566qnLLcMDK/S2226b3OJM1uaGNlxwLZl55pnLb0ErhJAOggYh3gyDffjhh+WWoSU37qzSZ5xxRpoIxU+ai8dw4V5MlBlqpAX/aJ2b+igKOhr8Dw3JD0ecWBOJNIrSJZh0Me9AJ1WUDtOIRFOIBXYmfdQb6u/hqsO5c7BAqyPkp+222y61KybcDxfyuvoyaJ0Q0kHQIIa/TBQh1oYD4kyEDhbgTgnBJUqFIfChhmuLoVGThrK/owbh+uuvL66++upixx13HJY00ijyGyeog0kXeZqvu1VR5aO55547ddCCSRvlU/2tHh8O5Ku77rorjZjBfA6T64erTQG/cXVW0DoRtSMIGoSQZlGwBPlQ+9+q+K+44orisssuS24DLGXcCIYT6cHC4zPDDDOUW4cGQtrzE9FWEmTlyYvlCMVnZczhQFpomITWiqgdkx7enzzFJ5rYYTUUj9xI1NixY9MksVjVdNKFkPaOuaQNxxwKoTGF6TSaZi0AE6KJ2GWXXXbYIkGprz7xiU9E3PsBEBbpIGiQ3q4dhKQKkR+lynkwYfkVvN8QMyGt8htq8j0QrZnerh2+W4LXBMjBRgQFMcefeOKJtDKX6B3C35kBPxR45yKovPzyyylt0Nu1w3fCTGSVoPPJZZpbxyyzzJI6sHlymPwm/m8w6UCkKp/Z4qrM1rt2qNNzGR4KdywCfrHFFktuZ9w5uOottNBCQ9Y5Y/l+6623UvQpzw55fDh9tEcCsbJhEDSIipZg404gZrOwbypDovHkk09OcbFHMibxXXTRRcWvfvWrZBEnLljoL7300mLfffdNQ+E6FSYAcq0Y7Aks3gfrDnG/yiqrjIvc4T5tH+zVJ4lnFqXTTjutWGGFFdKiONwAjBxYNY3F/Omnn077aChjGfUgGFpEXBED3CRxgpUbhfpJ2fU91+FEpdV0R/oiSgxBN954Y6qTlllmmeSyxEpu9GXvvfcu9wqaJYR0EDSIypcwYl0kJi1J/cILL6SZ/DvssEO5V3N85jOfKVZbbbXy29DAAqFD0CysGVZVNMRt4YBVV101DXuz7pj0d+uttxb33XdfEpOHH3546nBMCFZ1i++0CsuSBlHjZwZ+fYQO74m/9ECXmSfIPdOEUHWy7BxwwAFp4Q4hCJdYYonkdiI9WMotMf2Xv/yl2HLLLYv555+/PDJoJ6IODFf4x3Yg+gz3pKD9GC376U9/msop4Uw8EtMMAL/+9a9T+VafsxBvs8025VH9M+WUU6ay3gmwJj/44IPlt4mjDrcvg4hITzr8c8wxR6q/jO4FrRFCOggahEDjh2uyCIFERKuYWF5bDbXG3/qoo45K/yuKhhmJXEJzvfXWS9uh4mc90Qh861vfKre2hqFrIfOaxfMbAjXhka+oCphl2qQ/acEKrFK3qt8PfvCD5Hc3IfgDHnbYYel/IaAICbFUWY7AQsTSf8stt6S0INpNzGGFZkHS+HHl0FD6HcQzy4p7834GOlzq+joEE0NaXn755Wk0wnuxqqJ0MQtep4MfpA6FBny4Q26NVKS7EREoj0ZG5NX6UHXymI4Nlw1lTr5lfXz77beLhx56KOUhIwrf/e530/6Oz7/p7Bp94Xtfv52PbTs6wc5ndc6g/ejke1fc0dQ5CyywQCqjjAnqHJ1xdYo6fNFFFy2P6h9uPzvttFP5rVZXyHcEeZ4b4ZpWwlQ38D/m0sHVSx60FoB60mRW+WsgqJPPPPPM8tvEcX11knrSdT2HcqJTsO6665Z7Bc0SQjoIGkSFq2KERphFmoVahTh69OiJCscJwXLJoqaC46Ig4oRzmuR0wgknpH0UURaVXXbZpdh6660HvEQxkUoANgsL7fnnn5+sOJbeXn755ZPPNuEvxq6/LNIELXeHiS31np+bwBkzZkwK53fcccclwQxWXAvOiJWtwnctFb3GShppjIj2zTffvNhoo41SR8O+rE8aLpP9jBIMZAJP9qecEH7XubEgDBGmUdRQE/oaVMPKxLTRiw022KBYa621yiODduJ9E8dENIFiKN/7lwfhPRGrrHB8UpVXMXy53tjGp1+eJciNLhhR8d6vvfba1GlU1rnucBXi7z5q1Kg0HC4m8VZbbTXg2NLK/nBEvukGdLiPPfbY1AEilLnkmV+iLpNn1GXihBthO/LII9M7bQR5J68mK99dd911ycXtnHPOSfWe81vMx3b7Go3aYostkhVcfcfwIJ+p73Kd1yrNRN1Qr15zzTXFxRdfnOoo+Vo66FDstttu5V5B0xDSQRD0T1WsVaoNdaUqlNL3agVaueeeeyqnnnpqpVpRp22tUBW2lWoDXamK5PSpNvrlLzU++uijSrXBr1Qrvsr1119fbv041Qa5Um3g0/9V8VCpVq6VaoWevreDqtioVCvhdA/O7RrvvPNOpVopp9+lQVWUVKoCuFJtwNK2/nj//fcrO+64Y2Wuueaq3HjjjWmb53jmmWcqq6yySuUPf/hDpdroVNZbb72URlWxXHn++efTvVx44YWVqnCtVMV4pSqQKjvttFPllltuSWlw8MEHp3vtC+ktTaviJX13vWrHIr3fZqg2YOnezjzzzHHvzDmrQr/y29/+NqWP+89pFgwu0l6eqHZoKjvvvHO5tVKpiuJUfuSJN954o9xaqVQ7YpWq+En5tip6Kssuu2wqz96rfLbNNttU7rrrrnLvSqXakU75S15U9u+8886U5+TFvnBe15av5AX7VYVM+WswFKgzqp3/ypNPPpneh/rQu3300UfT7+qxame3Uu2Ap3qkFX75y1+mfFDt7Fd+97vfpW3VDnZlu+22q9x0003j8od84Ls6Xr3gurvsskuqe/rC/bo/dRXkvwnt2yiOr3YeKmPHjk33AGXC96B1IvxdEDQISy5LFdcBPnIsYSyyrLOs0a1YpMGiYKjNCldcRFgNWM24MrBWcWEwOYQF1/X6cllwb4YSTSRhHWUl4d7A0sVKV63Mk9vIQFZlZK1xbcOg3BWq9UeyBLNus6DzDWYB5qLByuF7f7A2m/Bi2N1f5zHs6p6lJxcR6SwNpLshSGnvXlgKL7nkkmSR9mwsPSJ2ZFcPFvK+rD3uuSrGk5XfkKs0Ysn2bqWzdGcpF6VhYrCqTzHFFOn9ezfwvvi8Smf34VzSi8tAI+kRtI78warsHZhUxf8TrHUsy6zSLJTyj4/3ww3He/ExPM/KKE8YHWKpNOKQ8332ZZ5tttnSO2fpNrmWNbOvUGqs35awl6eVT+fiGibyB4ulfOc+gsFDHaFe4VblHcsbyrY6Rdqrx7w/i1rlfNAM3iHXCnnDOzVqoU5TF/NFZulVv8uX6mCjZuoV4e7cCwu1OsLvvVGnGd1yj55D3jUKaoTLR/3oWo1a0aGMyN9clVwX7kuaSIegNaJm74XMrVE1dNzpEDJEDAGhIHQK1Z50GtLWyAwXKi/+tVwRxIQ1FDtQNJwqPpVkPa1UwPUQvSpdbgEqZcNuIj/k3/j49TeZiji0n+PlCxW7lQ+5iVikRFqcddZZ5d6tU/+crkOkGKasRwWvoWoV+YfbRq7YXZPokfYZwkRZJYQ0TMoBYWu41P4aH+K7L9yzNCGcnYMLhmFZMbp1aC688MKGw5z1fu/egwZPo5oZaHoEA0OeMNmTT7734/3qrNUjLxuC5zMq73DX4Bqi46azJi9x7SJusughYAiZvlaFU/8oi+ZTOK/656qrrkr5i7iW/5TzYHBR9urLqPei/u5dh7dSRp1LKDl1lTkQGXWTzhMXI/Nc7r777lS/y3PqnjwPRL5wzb7yj3PwZWYYUa+p3xgXuBaa7M3tiFsSo0szeE7nq8e55dWgdbpCSMuUJkIRVX19VKx6jnlfvUAWjU4mi+jTTz89TXognOohEPh/eT4dAxa/jN8UbL9dcMEFqVJvF87NT9bkHxbW4YAQIyqJR/fC902FNFBUyGY3Z+tju1Ahy39mlfOx23nnnZMIJvSIPFZPluiJwarAWsZ/2jtQwWv4NfYsaCr2di+aolJm4eCPOtToYPCXbnaCjPJN1LBIm/yjA6rDx3dSo2QbcdTqM2kY+UhKl6Az8E6UWe9UWEZ5h/jJqC/U9967smJ/Iyo+IhmwbCtbzaDsyp/8cgkm15PniCjXYOHur0wH7SfnhXbU4d6xUQcGkHq8b517kw6XXnrplIdYoptBfc5w4Fyia8g/8hNfa6NdRkSMnsizA4VleiAjlUGXCGmWRFZJvTiCmmXAGveG+wguFoc777wz7Svjnn322ZNEqCqFzXBhX3hmvUwTHg499NAUfcBwEHJv16QtE7omdI5WcF1DqM32lNuJdCFIiUpWAWGNNJYDhZBWAfc35N8sOkUw+UP+M8xIBGvcdXYMH8qj3ierBItnPVkcEs+GMQkFHSfPrxJmRWMJYb1tJ1lIt7sSzkLGfUOe0mnUiYF3yULIqsT1w3vRGEgH797+LMJ9DbezSMr7XGd8CGkdZ5NupJWyYOiTFbMV3HseMg46jzzUX18fyFtEbnYFqUe+Inp1dnVKiZdsZLGNmJJXe2O7kZocIYIbEUu2Dq18rXwPdpz14OOwxqq/B1qHM1YYteY+RlNwufCd9dm7zxDT4tsTvOp2f+U3qIvUP33lH/W5iEQ6YvIqq7V2QNugfncN7hnOOVDco7owaJ2uENIggE499dQkHPfaa6+UAbNF+ogjjij3mnQgYlhYJuTiriH3nIbz+cwS0Z5fwfXsm266abHPPvsU66+/fhLa7cJ1RSgwRDpcqHj4umarAL9Zs/QHispTg2jmfjuRZkSu5a2JQJUkMccSzaVBRU3sqUxZqFlB6lEhE84aCc9OUBtSZv0iMnfdddf01+gFodkusmtHOztiIM5nnXXW5KNKEBMufFbFrJY+8rL04E9OkBAsGgKWYC4ZuYNZP9yacT6dEaKGxYeVxzHyio6MpcXNam/WApnxLnR46l07gs4gd7CU4+ybTNQQP+pEgqe3S4/95Td1qDxCVBvNU86UQ7/3HukhsHX05ANCXMdXfWQ/5VmkD/Ww0cDeLibB4OLdEKgDrcN12n2cT/0s3xgVFgGm/p3KH/KYThMNwlc71w+szPzy1XX1OK/745aXfaONWMqj8pP2VdvA/a/e3a1V1K+NurIFfdM1kw01+oZg/CWG+EMeeOCBSZCyqKnYiBeWVBnUNiKMKNHr1PA6RqOde7P5ex4GhAqW7xIRIHNq3GX+3tTvxxoiM7u+yp5IIBwILNZzhSifx/0TWvnazqPhF4Krr56t8xFZ4p3mkGQmgymsCqGCrJFgnSceFHrP6p5MVnMtDQzrH98+FYG4uZ4tW2jGjBkz7rsCTkywdrsf96vhUcFki6hrq8zs4/nzb+6VtZBLBoFG8Kg8nLMeDSGhlEMXqWjqj5ce3FVYMD1fuyyxzi/NvBfWy3ZB5BKPRkzkAxUzNw/uBnyjWV3FvZVmQqixntZDOLJYs3Rp6KW/c8lP8kgeIvRuhZFrx3AgspA2AmGosRU0Ovz+fOQf96/BkR7KAUEi/7Musxhyw8iuSvKefErQGEHSkeDC453rdOgk1peJnO+UO5Zj5/Td+eUVftL2dx/+KifNQtirM6T9QK1eQXPI9+oheV99xcdefUeUqBPUGd4NlwrixXYuVFz7dNLkKXURS5+OqNFK+UseNTyvDGkvtAfKkrLF4tx7aF+dqe5koVRPKJ+G9h2rrmJtVOblFT7Y4QY0dBC+6knvYiCuNeoahgp1s482U11yyCGHJPGrnpKH5B/awntWx2i7CGTte86LvTv89lf3aQfUUfKKfEObuHedf9vcgzpqICE+oc0h6pWBoDW6QkjLdHniUm8hjfy7TH7KKack/17CU2GzWAYfW8Ja5ibeVJAaaxZEAsCQC1+oLI6JUtfwm0p1ySWXTNfJaNBZKPbbb790TRW4ytk1FbD9998/fSfYXEMjoFGW0VXg3BVU8u5BpWwm+ISEtPNz7xAj0j0RIXmp1HohrdBb5to+xJqKnwXb/RBxxx9/fJqsQ8y7d+ckYj27e/FdAVepaNDGjh07bghT40akEOSsMiocjZ37VpkQ5izYOb3FT2ZhdG2VFVGSIWZVKjoFGkJCy7tUSTmHeyD49fpZfwyDtXOpaBUxATfQyqseFaLnZaWQxwg5eaAe+VaDLJ/WD8PJc9KJcPQeWT50HHQCpZv0U1GyZBPmGv524n341L+jZvBMLIKeWToQ0p6PaJFHTVpVPq1S6K+85916Pu/f8QSzBoeVUb6V79Zcc800DFqPBko+tZ908juh431KO+JaXnVtk4T6Kk/9oWzLI7kjHgwd6h11g860/KD880dmUdZpJxaUW1FevCd1HZc++S3nJWXEPup5Qhn2z50inVD5gtHBfnyu61Hfup48asREnUeYcxWyP+HEcqkONGwfq10OLd67+kre6G2gGQjynjpaG638q8e1i/KDfJDdeIhsHSdGIvWQ2NL1HSn3R1/o9JmvQaBbCMi9ytPOo81lvNAWDDQGNbQh2l55NWiR6svvKqqFKMUGrTZy5ZYeqqKvUm2AK9WMXakWgkq1Ua1UM3Ol2sinGKTVAlKpis3xvleFd6VaOabz2r8qflPcynPOOSedq1pgK1WxWl6hRjXjVm6++eZKVQCm46rioFIVqClGcVU0V6piIp1z9OjRKV5pVURUfvjDH6bjqgK7Uq18U6zcauGtnHTSSZVq4axUC1959vH56KOPKnvssUeKnWufqqhP8XmrArRy7733VkaNGpX2qzYilW233bZSFdHpu+tWOxDpuo5bbrnlKlWBUdl8883TdS+55JKPfa82FilOZ7XnnPZfcMEFK1WhnM5d7TSk56o2IpWzzjorxf+VTp6x2tBUqg1YpdpTr1SFXqXaUKX/+8L5Pc9WW22VvlfFUWXvvfeuVBupFM8Tv//979O9VCuz9L1dSJMbb7wxxf/sFP76179Wzj777BQbdaiRd73fE088sdzS2VSFVKXaQUmxqwcL5652dCdYHoORjbpPrOkrrrii3BJ0ElURmtr/22+/vdzSWWhj7rvvvhSbfqiodhhTOxy0Ttf4SDcCS1T2l2b90vsTNsl2k/X02lgW6r+zTrAK60kasmGFyj6thqg33njjZGmsh+Vr5ZVXThEHWD1YnfN2w9cs2CbEsHa4jzzxSe+W5dg+rBv278sPtC/cK59qQ0/ZX7oR/zzXdxyLtmdzvG2e23f+1fm7NGD9BAuj4SyWSpZ1K9+xFBqGl04s1dKJhZFbgOFR1iO+246d0DCT46wWVe0MpO8sRFUxn94JC8Bg4xmr5ab8NvzIA6z8rF5DjXTwkSaTAkZTlK1cngaDnCadlEeCoUNdyMKt7gs6k06rw3vDfdII91AxKdXhnUoI6TZDUOZJjPzvTOgznFOPTGv4kW8e948spPvDkJQhesK0FYguQ/vCq3GH4D4yVHCxIOYNqbkPw5o5nURJMXzaCAq9cxHl0HAZ9uLaYUhtMOF6YKhNRdcp6EiodIfDjcD7lLeHQ8S3gnvlIz6YKJvcU3qX+aA7UL/xW82TGYPOgpFG/d1JdXg93Dws3qQOGSoY/IYzOMBIIIR0myAq+BixuPL5BAuyiYu9LdK2C8dHSPPNPOOMM9J2Apvf3oQgGl0j+2Dbn58zHydWWj6g/cFyy0q+xhprJH/pjPsnxvK9ukfWYudvJYIBwZvvx/3xXWVl5ufFws0HzMQesDJLi0ZQEbLWm5CYRwL8zdsHk/xMfCmDGt4tv/2ghvxoXoR0CYKgs1A+1d9Rh/fAv5vfddA6XbVEuEJkNrUJJqzAJmIRYMQdkSQziUBhEQ8WBRNM8mxv+xoaZsnt67tJJKIpmKxkop3zmrFrYonJe/UQqYSvfbhomLQnsoVJT8Ql1wfHOaeoCM5H0BrCN0HKZDoTEkwUdKxncR5uHtky6XnMXBf1w8QG31nLfViEnYdV3DWE/QJXD8/jPohoq3ARSc7JEm5SpElUhsbdk5nJvuvR5u96+lw0HGfiH+uxezT5Rgg6EySc37nzZEW/OaftOh7SUIehr2gbOhPuR2eFVVo6mLTIDYf7iGcykdE7liaEb7t698SRyUzykXRrFu/dxECRJaSNdzEYkR00EiZwmuU9mBNI5CnvWV6xElyjeCfyv3wuf+d7zNvlIx1Slpl2Iz9yKXINEw11LNuJtJevPZP3GwwN3quyyRCgLlFWTWQWvUfdxdKXXXqUCy5y3lP99nZh5FB9bcIiwjrdOcgnXBsZb5qZIK3uNsGPyyZDkLa7Hm2xOoVbT+/fBoq60Mi1utaIaLsxUV27FBNfW6erhLQKjohRyZkJa+Y0QZwjerAkmd3tN6KSwJbBCDqiVDB9oiF/J2xVxr6bES5iBdcJYtg1FAB+zr0ratZfjaywW/ZzrOOIZ5EKFFp/7Uf0sj77roAKw6SwOlYBYOX1/dhjj03CMUPkODchbZjZNYhNwtd5iVZDkIaiVSjcFjT+GiPHuRcLmThGNBHRDgzha4Tsz8LsOyFc/11Dxg/VjGPXlF4EL5G77LLLjnPFcEx+fuc44IADUlrzGReaipW5rwUS3CeB5RwEtPcgLQ866KD0fglUkR6IecJMb9us6XYgTZ3T8K00bwbHeibvQ4Xr3r1XEVTaLea8I9FPvEvRKwYLz0SwEI/ySSNwv5EndAaVEx1IHUD5go878WG7URD5Sb5vJxpSdYCY2spSuzsy8qDOQe5oB0ODeuS4444bZyRQ53Ctk6dE5CCm1bHqVmJIh135s59h7XaFhIQ8oC6Tx/zvukFnwAhCRHvfjdbh3iEDzYknnpg6+trDetctdQqhaxEw4Urb7dZF+J955pnjomK1G/evXqZnghapNoZBEDSA6CSPPvpopSqCyy2NU62MK9XGvlIV0in6ysMPP1ypdthSxJZ2U20oUnSXTTbZpNwyOHimameuMnbs2HJL/1Q7WpWqiE7RLaqdoBTZptqhStFHpI3tIrvstttuKYrMYCDSyBJLLJHeR7vxHNJehJBgaJCnLr/88hQp6KKLLkrbnn322Uq1A12pipDKc889V1lqqaVSpCLRVHbffffKnXfemd7/oYcemiIotRt5WPSW448/vtwSdAJ/+9vfUkSoJ598stzSP+p99fXyyy9fWXTRRVOdV488ttNOO6Xfe//WDv7+97+n/L3FFluUW9rL22+/Xal2EMpvQSt0lUU6CAaCXjs3GqMVzU7OMArA+snant1TuP6wrucRkQyLCdcU1jSWNEPDfMKNfrCocaXxO5cioyT+clligWadZwk1DMllhkU6n49vvVEClgeWdVY5VnIjAq1Yfll3jIqwIhttaAQjCkZ6pAVroDQ18dR9SxuWIvv4cP+xilc9LOCsfSbKel5pafTEd0P5hl2NUrAQGcGxv1EAox+e2dCokSdD/izS3oPzWOJXTHJWKteW1tLf/Ti/yayNYDTAuzDi0ugxQetkFw7uOsqC0SIWaUPt8qXRDu4b3rFIGkYJWRWNFNrXiJXRtt6TUA2jG7ngziY/Ge3zndtZtd1M5+QewlJplE9e4RLIeih/w8iK87NIi2YkjyqryiMXOPnfvSiDeQQ0GFzUAd6hOqD3ioITQn1ghEk9zE1ynXXWGWd1VneqW7xD57ZmQW+LtH3kD/lMXjICaURSnjWCqz733WisetFISa6P1G/qRu2AfM4i7Rijmtwb5XN5KbsrqRvVWTmPNoLruL+INNM6MdkwCBokV6gazoFCWGvIe/sBEwZcH/icqxhHjRqVKk2NtEVa/G8oTqNM1Kt0+fUTnRYD4h9ej/MRhfZ3PsOPBLZG3oRX2w1ZtkJ+hmaidkhDxxAoIrYQqb2j0GgEDNH3DoGYhbvjPC9/fv9LA0v/W0yJILHPlVdemRof+xDVRNXRRx893iQj59Ox0KFwPn+5dmmUpA33Er7mGs9G8SxZ0AWDDzcaQ95cpOoheggD4Uy9P//rLBJQOljEizzmQ6DUQxARPcqS8mHxJ3lJHrIoFcHjPDq33ER0iJVXHSj50bZ6CB8uTI73Mcnb3A7HyZ/m4VhkKxh8iFj5oB1ROxgB5B11yIQMCepq9bnOvPzi3cuPRLT6ihuiOkl9qA5SL5t47391kDq9HtfUKeQaJ79Z0da5CGh5yXbHqAMbJaJ2DJwQ0kHQIIQja2+e0NkqrMosEyrz3pMWVaqspSaoEr0sZywM4pYLc8cyRgjwQbfiJmHNikFI8jO3bz3Z8kwwmFSqYldBs1izyJhgMpBGRcPU7GQtz29+gnsgQAiTeljsWElElqlHI0I0EU8Ei5jmGkXpopPhObwbnZ0ddtghdVI0SGeddVZatZPgZyHMOB8LIdHEKk58XXDBBckaqXEU31zaEsaNoqPAgtTuCUfBx/Eu+T8rl707c0YDWAd1sviXNjNx1bsncMy7GD169DgLpPKl3BEe6gHnVz6VQduF8dx6663T/dRD1CiDyroyR/QQQa7jvnUY2z0XIOibPBrYjvkLLM1GOCY2Sc+ogw4Toa0e2mSTTVI9tfnmm6d1JOQldYW6eaeddkqdLh/1+d577/2xiao6cKzH8o4J3uownX3ths67fJit2I2i89/M/sHHCSEdBA1i0olJTURwq7C2ssJys+jttgAWZMPD3C9U9uJrW6JdQ+5/DTJxrAIlSDXSGmeC1qRKDXk9zseCwQLGMmJCKfcG7iSst4YGCcZW8CxErYaiGTRkxInJWBoQQ6MZIpq49byG6OvxLIZQiQ+NjwZMY2MI08RZacCy43yeU0MnDQl9Lhsmo9WLfucjxDwDK6JOBsulTofzSS+CrJmJpcQdq5LGMBhcdHgMgeuUEROGx4laQ/fKmJEYHVCdJB0kokd+UI7lfeWHAOm9VLR8QKgQvgSuMmXysv+5gLD65TJoX3mSUCdGVl999Y9NknYtHUAfHUST0wkk5VA+kf965/VgcPDO1N/yzECQdxgC5D8jg6zN6lijWOqdjPxlhEteYgThmsHdSJ3incsT6nv3JP/IVzru6jL5dvfddy/PVMP51Fn2Z4CQn+XN7JKmfRIGthljj3JklDJonRDSQdAgLE0E3kCG7TWqLM4qVZYJIeDqyRbNLC6zEFaxiiaj0mVB9b993Q/Bl/dl7arHPkSlqCnEhGFqsctZQrbffvtUAbPYER7NIj3cV28h0igEMBGfxW22EPsQLISPRiPjWVjcc5rZ35A7RKHRQBmO15DxUWZp0VHgn0o85f8zzufeCXOinsWIpcj7lUYskEQTd49GcU7PI12CwYXlDYSzqEGEDHHDCu2vvKBzydJHgCgb8ruyR8AQOLb1juqjkyaf2QfKrCF8+YLIIYaVOcPh9pXPeu9bj7xgX9ZrZZC7iVET/vxbbLFFKgeG8wmaYHBRPr3HgdTh4BamTtHx57bDmKAOJUjltYy8IZ/melnHSf6UJ9TLOuo6/+p8+7o/dZoOmrxE8Ps/Yx8dOtFB5CUjbf5Xn1sfgqjm1pbzYyPIfzGfY2DEZMMOgoWPCOBPxQ+3HcNPA0WFofdrog1xMtQCwfVVJnr8evXDKVC8H0NrevvNWCnhOVgL+LQRswQki5kKuL4hJ04JYuJNpcvqIE+oIPP1WU+JYBW086o4swg1+Ymli/uGypvVg7AbM2ZMsqK4HiHAisbtQcWswuZjqjJuBvejIXFPjYa/08joSGg8CCCNBAHsvfJHJSjcJ8FrCJPgyGnteTVe0sZf6cf6a4iTFVnasUyyCLK421+a6IgQVtLShC4WJH7TGiQdEuWNVdC5NITENet1bnRdq9GJOPnedZI6ofyOZLwbZYeVj/VO2ssLJpHqhMljxI1yII+K869eVb68f1ZnZYsbFReejHxEZPNndrz8Iw+o/5Q351bONt1005TH5B2WSX/laWVL3pFP5QUWaMcT9iyOOslGknSK5UV5V1laYIEFxruPoP3II96B+qaZOtz7Uqeqc8SftzaB/CDv+RDF2qlDDz10vDk08oE8ZLK3POjdqwMd7x507tVzRieJWb/lNRLs65yErryko6g+lz/Vlep8ozDykXr40ksvTR1A+cm9uadGcE2fCH/XOiGkG0RFp+LV6GarmUZXQ6xiJlTydgVAQ96K6FPoiC3D1vXD0MOBZ9YQnHDCCWmiloZjQr5UGgoiTQOV04a1VEOl8mpFVLi+Run4449PwoZ/2YSuPxR4zxpKFZiKqhmkj4pQBUjoEtXSVuNe7yetEmSpkoYacJUvYUDkqkD9znLF3UMjbrv0NeHE+QgKQt/EQkLREDL/PFYO5yMQNtxww2RJk9dYLljZxEZtlvx+uKksvPDC5daJo3NA7BI3hIdnI8JV5PxSbeMeoQFxj6wsGc8rT7E+G0L1vPxLHe836cMayHdVPlH+NGr21RDaRnjpQOQhflFNiBeCRroqd9w6vGMdFsJp/fXX/5iv4oTQSEsP73g482q34V16Z943AaFcqD+N3ngn3nuO4GE7C7a8RgT19q9WfnS4TPBVTp1bPiVS5DMQLvK8POZaRk7Uf/IuP9XcCXYt1mgjHPKT88mn/GOdl5BSL+goNxr5JmgdHXeGBHmid7SkieG9qUeUa+JYvSMvZbx3dUXv7f5XXxG7eS6IdRaMivjNce5nvfXWS7/pHMpnxLX8SXDr2Puuc+5/+U7+48YEnXznk5fU88rAKqusMt59TAx5V3vTqotfUO18VxvDSvl/MBEUEhYrgk5DTKQoNCaYKAz86FhAFFQNuQUxZO5OhSgkvhTqCSFrGIayMIueb+6N90YDpscslFP2zVLZ8N1VAWmsCL9mkeYaGSsiKuiG9BvtZQ8G3nO24rbyPAPF9Qk+wo/YG268H+/XaMXOO+9cbh0+CGERELbaaqtyy9Cj48PibgKkRjcYWRA36kF1O/EbTFp4f9xy1F3K6HCi3TSyoZPPPWO4YPTS+e89vyZonPCRbhCWCBWnSAqs0IZiiGgQVlbRIkqJa6GMOllEs4RoDMxInxgsJ4bWe094qMe5iOy99toriWhD8z5nnHFGsh7miRStIM2JkV133bXcMrzoHDQzZNYudHpU/kYqdOY6QURD/iDqWduGE42jsFLcf4Z7eJIVyFA+K1QwcuD+xIo9duzY1HkMET1pYgRBmzKcBhkCmni9+OKL0+h1o/GsBwtaxQTFoHVCSA8ier2G+zTyPoRQxnC84Xc9wfyb4UCi0/+GnojU/Hv9hy8UCCyWYNsUyjzUw5LMOuc83FGEWhozZkwaqnRdkyO4SxC59uGPZf98fucijhtBAyMOsWFsLiAZnQsTaY455pjk++UenNv1NETZHcF34tB3Vmf7iIPJBWJC2FdHIN+r4dv67c7JBaP3RL6B4n1wOZCmQ4nrssx7J436Ig8F8pk828zElsHAKJA8oFFq1Jd5sDBqwMqk/AYjh2w9VFc14xIQdBbaTD7urMDDhXvI7hRc9bhsDCfcL7n9Ba0Trh1NwjeJXyW/uPrVsIg4AdFZokwqIaJVvMQlIZSFoxnbfC6J2V122SX54rH66invscceybLNok0Imgxx8MEHJ19W5+P/ySoivm5eaIJVXI+SoHFvXN5ZzLmgELHOqXF3LB8qE9NMjDHb1/4mZrH48t866aSTkk8WocvSSJCysPFdFXqtt2uHrGNfxxgWEvmgLwgd1yN6WandM4uOaBGGwUVHILZN5uDDq9EiGk3Q4ELjOTfffPMkjFU6OieEufRVKXE/kW7eybHHHptEjPtUUfFpbxfSS1pIk94roXUj8rW015nbZ599yq3dDb9tZay373sQBMMP0cjgpO7ighkUqe1niOgE97xJlbBItwBRa4KAzJc/Viuqt1QSzoKqE4VcHSwgQUDz92VdJAJZgRVsvxOXJhnkCQnQW81hblh984QUE/8IWKtsEcGO9zvLMqHu2kSnykJPc7vttksWaBY7PWETuLihmFgl5Bd3BfdpgQ/36Zyeh4CfGNKBcODyMLFFKzzXnnvumZ6dEM4TNsxAJvQXXnjh1HkwMSenBf+1vq5PlBPgLEOsjzn6BRHOysAFQrpIq3b39N2zex9uC0KnwLVDx4grQ1DDSIxRA+nSTejIG/FSL/bGb9xudGqNuOXveQRMRyy7f6lPbDPqxmjQG/WlkTwjYUHQLAxW6m8TuoMaDFCxsuHACCHdAgQuH2miL39YROvDmLGUWjxDgH6IQGDSHlHJXYOYZTnOxxAlCjjBmXEdlk/nYoHWkyaUWbpYZYlxQjsfy2pLABPQxKRG3YIVFguYmM+2ysX9mECn8aoX8xPDdUU/YJkWdWFiuIbIEDoAJux5JpMzF1lkkSTiNcKseCBCCHz+5r2xL2u+hlcHhogWhcJM5RyqjCjX0AoR1050HHLnJ6jBSt+qD/xIRCfW0LF06RYIY2JY6C+jbvUoL+pH7lrqFp1j6UMMK79GeNRtOvnqEJERdOYJbX/rh+DzZFt1oEmdQdAs2gf1d+SfHrSVQ+2uONIIIT2IyKCsxCA6ha7x0SA0ioIv9A1xaPicFZlwdQ5/hR+DiXk5JFuzjbhrcIPgR61ha9S32DWFBeNGIbRTb79Q96fS4qZhX2LfwiDZT1rngsC3H0tzo1YmrhVbbrnluE4MC7X4sSaQmPTI3UAjzK3GddpFCOnx8d5CSI9PFtLNlPFJHWVX2C3PXg+BLaKLeMxCVyqPRop0lHfbbbdUdk899dQ0xK5uyLHN1XNGxxgC8rwPcPvS4e6mtA3aizyq/o46vAcd2BDSAyOE9CBBOHI74I+sgSA6iGrbG426QLixuPJ11thwDSF6uS/kgO5cGvK+3Dacu7+IIfWWZBEPNIKjRo1Kvp2rrrpq8rOGc5qQODFY2K0cxp9Zw5jFtHMbpmWVtxgG3C8LO/9vHQPuGyCo3bcGN8Ni3Zeg517Bp5zlSrq6RxMATU5UIXAPIaL333//ZLWXVu3CCIFOQx4WzNdmIfdeug35iC99zPjuQSfPLPxucu0wz2OHHXZIC4pklA3zMtRPyrZ6QblXhsz9yKEBiWLlWCxn+clx6g37Kcu5LlO2TWq1zWdCKIc6dgQ5XFcnn/Wb1Vxd5z6C7kTnTP2tDelGGKvE8OcaaXQX5ieFe97AiAVZGoQw1Gvj52dYktBjjeOeoZebo2IQy0Sqmd0yKIFpOJMgVaFzsyCIbTcpUWbmX8w1QQOQfQMVdr5LXg/RyEVEI0AYWtBCrFznJX5dj2gkWFl+HKcB4+bhvK7pvglV3/lDOVZjo+H3cT/umahVyDyjfbPbBTcMlQ+LEkGc0eA5n0bTBEDp4j7dDyu39LA0LnQiTMbkR0kkm0iZt7sHaaiic5yhXhYoQi27tbi+Btc5CHS/S1cVg/egEdXpcA8aY1iEwYTFdpAbaXlBgy993YdGmu+6fCC9uuVDBLHs8PnnbtTXPt32IdyUQ2JPWeprn5Hykd89I3TIuawpazpWrNTqDNsIbfWWkSmLleh8w/E6oj5GlNQDhtzHjh2b/lcXrLPOOmm//7+9e3eRotvCOFwnFQNDjcXMRBC8MAYKigiCMiAaeAvETAQFEzEY8IagIEZe8IqIkaiBgggiiAgiCCYGmir+A2bn8OxyO21/zUfbM3pmut4fNI7T1TU9PbV3vXvtd61lfjEvGM/mKvPhoBKDhIL50lynKYXdqePHj5c5jU3EHM4SJy+DOB/0e+Uxvg9/c0n3vjZG+58f94dFq+CeMWaMGmful/SA4FwYjVTtGBLCyWTcX+JNZJWgltBXITQlBBK0IqUEs2gLcczf54K2pSnCIsJKhOls5P+SBuEGtXfv3pKw2IvzEJRTU1Pl57pJGASOd9PhmRaZPnHiRDneexQxVpEDBKsEP6+9cOFCiQw5h8GloYrzWwA4p2NFmlTcgBug9z8o4k1UEe+is3AeVov+dZrjRIbcMKvAhvfj9WwsENHzGYke+Rc80M7n33osIa+OsURGN2QLEQmW9fuz6ZM28ViQ+DkWCP62hDwRoKpJ1zAmaotb115o7QwWWK69320jP98wT7BqwZgwd4k+m7csZI1RwtUYJHCNd3NN3YmyCNMO2VivVXAsylQP8HpBAfOP41xjtWIQ64ecFHaQfrwPycoscFu2bCmvc7yFNhFv/jF/2i3UvCd0C0Ja4MXc5RrpGq5/C1z3STZTeVECaAS1e3sYjQjp8FdxQ9WsRcvd+VaP1QLIQkFkTZSeyCckVWmoiZJdwtRhYiZ6BomaLiJ6ahGqrrqF6Dhjx8qiHP1C2mcgF0JQgZAWDZbLQNBqj426wyfRWdDBIsTujnOJ7EtctHAWbLh48WJJTLYjZBeIx1rH1F6bR7W9KYHpZxEHdrNcn0SDBfaqVavKe7TTxc4WuoXx6doyd7nmuoZ7mICgXRtzFEuHXV62LOM2jEaEdPjjuMHZmpVxLxJge2k+1h22BcZy4gYtOq8GNmHtJm1nQhS8S/hbEkwWFqJ/ofXkivi4QbkuukK/kBb5k7is+gbB6jpRZ14Em5h17bBYiArLZ4BIoZ00D9HuuhvHolFFr50stjALcYnF1WsNn70x6UHEE9UE9eTkZIl6E/4W8cR93fkL3UIgx66H66+LvuBqnRKRtjA1b9s5Y4GyMx5GI8mG4Y9jrSYixZPN66zj4XzEgoCVQySNr100zg1ZCUPPdQ1/V95YfvjQIkIv4iO62hWIE+Pa7028WjTL2xB9lsdw+fLlIm6NkVpvnk1KdLl3J2PBggUlwqyOtNwPFXf4rYnzWnP65MmT5bzHjh37RUTDtSi/RGUdfmqv937sHBHQLDe8/KKSoZuIyFr0eXQRQSDJ0MaRcpUTExNl0StAFEYnyYbhj2Pw8jfqyCi65IY5HxHFsE1MJPC7+71EztzsuxaNrhBEPhPNdUK7a8E/T7B1pXKHRYPdJkLWTg2B61HHicQ/n8u+fftK3gT83+skL7NZwPH8y7adLVZ9rfZ+L4QQ4c7jXJMW4XwWuYSznQBlOSVBi8BJdpRIRegT9vz8/SI8dAOLKNed3CHXV9dgNzMGXf/1nuXzsJvD4hFGI9aOEIbEJMxnKbEzGc7TJQ5FpFVTCG0yk2goEfdvZdrC7MI6ImHaAqa3MVYIvVj426kwd8ltCU3ZLVZJK+NmdGLtCGFICGleMlVRwrS1g3AMLawdqu/4XMLfw7XI+5x6uOHfqNaO2WzUNd8RDIm1Y2ZESIcwJEr62Q5TRSC0sLf01hXvOq4ROxY+l/D3YOfYtWtXJysxhOExPs3fXbXiDcJcVevBh9HIbB/CkJiAtWGvPs+u46bE36pmcmjhQRQVHdQsJITw/8Wi3/ydOXwafSHSnXZmREiHMCSqDtgWlAgV2u10SSqSuEILa4eybj6XcUbirbFw69atUqtZtQxI5tNwSfm52qYbbFF8mI5XO1plj9nGZ69ChwZYfJ8h9CMp1fydOXwaDY+UngyjEyEdwpBU4SihLLSfB88hj11osdhyY3LDHmdUziCedSbUnEgSrnGhicrTp09LuTudUwlbuEZu3rxZytp5Tt1155hNiPUPHz6UetXxfIZBGJ+u03Ff6P4OFqBKRobRiZAOYUhYO5QNShe/FtYOJd6S4DWNslqqAYxz6TvRaMlaBLNSckSxJixuyB5nz54tIlrJy+vXr5fXKAkoQn3p0qXSjIkIn+2ooPJ5a9euLV3aQhgEa4f5W1nG0CKvQG3pMDoR0iEMCQFh5S7iGFoIp2yjTyMq+uXLl+b79+8/vjN++B2NAfVnr1271jx8+LBEl5X72759e7kxe2zYsOGnWLbogteo/6wxS3/CV69d5N69e82rV69+2kFEsZW4UzHn/v37JeLsPbCReF7pu35EHx3vecd9+vTpF/sHC44IdugOdccoc/g0xq45K4xOhHQIQ1KFtCYPobV2qMva1S5hg6hCmmAbV2T5q5NNRO/evbsIVW3i+5F4WRv1aIpCWE9NTZUOg+vWrftHwpexRUA/evSoCN8zZ84U//2VK1eaU6dOFf+1boiOIYBfvHhRRDVRfP78+X8s6JzP8+wnDx48KB0WXau+p3259uSDBHgYX+oiMHP4NKwuCYbMjHQ2DGFIaukkXdPSbKP9PIiqhQsXJgu+B/YOW8e9nffGCX9zv5uSWf7uKrcQtYRyhVjRNnz9+vVlvPhMXCd3794tXRD379//i0XKIlXCE5FM8GoOIZoswi16/fnz52ZycrJ0RfUzdUS8fft2c/To0WbHjh1lXCqB5+f4uWwlBMK5c+dKWTzvmeDWXlz3wzVr1pTXLFu27Gfb8jD+mLNctypV6Eob2s9ElaEudnqcLSKkQxgSN2M364joFhMwQRURPY2bNIE4riK6H78v3ylxvGnTpvI9Avbdu3cl+lfF9bdv35pnz54VMcz2Quwqm1i95JJWWS0kLe7cubNZtGhR6Zbpeef/+PFjeZ0kTsLcv6LMBw4cKDaSlStXlqi3qLVzW8jYLVEhxM6JCKQSX/z8rtv37983S5cuLZF1rwvdgJ3I/B0RPY0FbkT0zIi1I4QQwkjwV4oWE7IgdnW61N1RNJrNRWRZR1CiVqT58OHDRWzXih4QHSaYJSWyZBDh9WuiZ/Xq1aXix9evX5vly5eXY0Wn/RwQzb0l9ZxPlM2xp0+fbq5evdocOXKkWbx4cUlGPHToUEl4vHHjxo9XhBDCaCQiHUIIYWiIZxFodg6imVjetm1bEb+PHz9u7ty5U5K6JAe+efOmiFfWjdevXxfLh8izCLUItugy7PY4xvk8TxQTyXY77AJ5jm9648aNJZIsquxcT548KdFmkWxt2ZXZ8x5EylUi4KUm2HmrJSjyrqt77f2JxBHqmzdvLu8hhBBGIRHpEEIIQyPqzBrBqkHsShxkrxAV5nMWDRY5fvnyZRG3K1asKJ7mgwcPNm/fvi3iVrS6v2zikiVLSvIiG4d61M6n3CT4sIlox0CUeuvWreWY+j6cj3j3nJ/LFqIsH6HvfOwgExMTJXpOVIuSK98XQggz4T//ZSALIYQQ5ijEsEobe/bs+fGdEEKYG0RIhxBCmJOwbzx//rzYSSQF1oTGEEKYK8TaEUIIYU6ilTMvNutGOhaGEOYiiUiHEEIIIYQwAolIhxBCCCGEMAIR0iGEEEIIIfw2TfM/ecMSSXKlsDoAAAAASUVORK5CYII=
*/
